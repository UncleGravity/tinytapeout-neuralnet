/*
 * Layer 1 Full - Complete first layer with integrated ROM
 * 
 * Self-contained module that processes all 48 neurons sequentially.
 * Weights and biases are stored in internal ROM (loaded from hex files).
 * 
 * Input: 64-pixel array reference (no cyclical management needed)
 * Output: 48 activated values stored internally, readable after done
 * 
 * Architecture:
 *   - Internal ROM: W1 weights (3,072 entries) + b1 biases (48 entries)
 *   - Reuses 1 layer1_neuron module for all 48 neurons
 *   - Reuses 1 sign_activation module
 *   - FSM manages sequential processing and ROM addressing
 *   - Reads pixels directly from input array using mac_count as index
 * 
 * Memory:
 *   - W1: 3,072 weights × 2 bits = 6,144 bits
 *   - b1: 48 biases × 4 bits = 192 bits
 *   - Output buffer: 48 × 2 bits = 96 bits
 *   - Total: 6,432 bits (804 bytes)
 * 
 * Timing:
 *   - Each neuron: ~67 cycles (64 MACs + bias + overhead)
 *   - Total: ~3,216 cycles for all 48 neurons
 */

module layer1_full (
    input  wire        clk,
    input  wire        rst_n,
    input  wire        start,              // Start layer 1 computation
    input  wire [127:0] pixels_flat,       // Input pixels as flat vector (64 × 2-bit = 128 bits)
    output reg         done,               // Computation complete
    output reg         busy,               // Currently computing
    // Read interface for outputs (after done=1)
    input  wire [5:0]  read_addr,          // Which output to read (0-47)
    output wire signed [1:0] read_data     // Output value at read_addr
);

    // ========================================================================
    // Unpack flat pixel vector into array
    // ========================================================================
    reg [1:0] pixels [0:63];
    integer k;
    always @(*) begin
        for (k = 0; k < 64; k = k + 1) begin
            pixels[k] = pixels_flat[k*2 +: 2];
        end
    end

    // ========================================================================
    // Weight and Bias ROM
    // ========================================================================
    
    // Layer 1 Weight ROM: 3,072 weights (48 neurons × 64 inputs)
    // Column-major: neuron N weights at addresses [N*64, N*64+63]
    reg [1:0] w1_rom [0:3071];
    
    // Layer 1 Bias ROM: 48 biases
    reg [3:0] b1_rom [0:47];
    
    // Inline initialization - generated from weights.npz
    // This works for both RTL and gate-level simulation
    initial begin
        // Weights (3,072 entries: 48 neurons × 64 inputs)
        // Weights    0-  15
        w1_rom[   0] = 2'b00;
        w1_rom[   1] = 2'b00;
        w1_rom[   2] = 2'b00;
        w1_rom[   3] = 2'b00;
        w1_rom[   4] = 2'b00;
        w1_rom[   5] = 2'b00;
        w1_rom[   6] = 2'b00;
        w1_rom[   7] = 2'b01;
        w1_rom[   8] = 2'b11;
        w1_rom[   9] = 2'b00;
        w1_rom[  10] = 2'b00;
        w1_rom[  11] = 2'b00;
        w1_rom[  12] = 2'b11;
        w1_rom[  13] = 2'b00;
        w1_rom[  14] = 2'b00;
        w1_rom[  15] = 2'b01;
        // Weights   16-  31
        w1_rom[  16] = 2'b00;
        w1_rom[  17] = 2'b01;
        w1_rom[  18] = 2'b00;
        w1_rom[  19] = 2'b11;
        w1_rom[  20] = 2'b11;
        w1_rom[  21] = 2'b00;
        w1_rom[  22] = 2'b01;
        w1_rom[  23] = 2'b01;
        w1_rom[  24] = 2'b11;
        w1_rom[  25] = 2'b11;
        w1_rom[  26] = 2'b11;
        w1_rom[  27] = 2'b11;
        w1_rom[  28] = 2'b00;
        w1_rom[  29] = 2'b00;
        w1_rom[  30] = 2'b11;
        w1_rom[  31] = 2'b01;
        // Weights   32-  47
        w1_rom[  32] = 2'b01;
        w1_rom[  33] = 2'b11;
        w1_rom[  34] = 2'b00;
        w1_rom[  35] = 2'b00;
        w1_rom[  36] = 2'b00;
        w1_rom[  37] = 2'b00;
        w1_rom[  38] = 2'b11;
        w1_rom[  39] = 2'b01;
        w1_rom[  40] = 2'b00;
        w1_rom[  41] = 2'b01;
        w1_rom[  42] = 2'b00;
        w1_rom[  43] = 2'b11;
        w1_rom[  44] = 2'b01;
        w1_rom[  45] = 2'b01;
        w1_rom[  46] = 2'b01;
        w1_rom[  47] = 2'b01;
        // Weights   48-  63
        w1_rom[  48] = 2'b00;
        w1_rom[  49] = 2'b01;
        w1_rom[  50] = 2'b01;
        w1_rom[  51] = 2'b00;
        w1_rom[  52] = 2'b00;
        w1_rom[  53] = 2'b01;
        w1_rom[  54] = 2'b01;
        w1_rom[  55] = 2'b01;
        w1_rom[  56] = 2'b11;
        w1_rom[  57] = 2'b00;
        w1_rom[  58] = 2'b11;
        w1_rom[  59] = 2'b00;
        w1_rom[  60] = 2'b11;
        w1_rom[  61] = 2'b11;
        w1_rom[  62] = 2'b11;
        w1_rom[  63] = 2'b00;
        // Weights   64-  79
        w1_rom[  64] = 2'b00;
        w1_rom[  65] = 2'b00;
        w1_rom[  66] = 2'b01;
        w1_rom[  67] = 2'b01;
        w1_rom[  68] = 2'b01;
        w1_rom[  69] = 2'b01;
        w1_rom[  70] = 2'b01;
        w1_rom[  71] = 2'b00;
        w1_rom[  72] = 2'b00;
        w1_rom[  73] = 2'b00;
        w1_rom[  74] = 2'b00;
        w1_rom[  75] = 2'b00;
        w1_rom[  76] = 2'b11;
        w1_rom[  77] = 2'b00;
        w1_rom[  78] = 2'b01;
        w1_rom[  79] = 2'b11;
        // Weights   80-  95
        w1_rom[  80] = 2'b00;
        w1_rom[  81] = 2'b11;
        w1_rom[  82] = 2'b00;
        w1_rom[  83] = 2'b00;
        w1_rom[  84] = 2'b00;
        w1_rom[  85] = 2'b11;
        w1_rom[  86] = 2'b11;
        w1_rom[  87] = 2'b00;
        w1_rom[  88] = 2'b00;
        w1_rom[  89] = 2'b01;
        w1_rom[  90] = 2'b00;
        w1_rom[  91] = 2'b00;
        w1_rom[  92] = 2'b01;
        w1_rom[  93] = 2'b11;
        w1_rom[  94] = 2'b00;
        w1_rom[  95] = 2'b00;
        // Weights   96- 111
        w1_rom[  96] = 2'b11;
        w1_rom[  97] = 2'b11;
        w1_rom[  98] = 2'b11;
        w1_rom[  99] = 2'b00;
        w1_rom[ 100] = 2'b01;
        w1_rom[ 101] = 2'b11;
        w1_rom[ 102] = 2'b00;
        w1_rom[ 103] = 2'b00;
        w1_rom[ 104] = 2'b00;
        w1_rom[ 105] = 2'b11;
        w1_rom[ 106] = 2'b00;
        w1_rom[ 107] = 2'b01;
        w1_rom[ 108] = 2'b00;
        w1_rom[ 109] = 2'b11;
        w1_rom[ 110] = 2'b00;
        w1_rom[ 111] = 2'b11;
        // Weights  112- 127
        w1_rom[ 112] = 2'b00;
        w1_rom[ 113] = 2'b00;
        w1_rom[ 114] = 2'b01;
        w1_rom[ 115] = 2'b00;
        w1_rom[ 116] = 2'b00;
        w1_rom[ 117] = 2'b00;
        w1_rom[ 118] = 2'b00;
        w1_rom[ 119] = 2'b01;
        w1_rom[ 120] = 2'b11;
        w1_rom[ 121] = 2'b11;
        w1_rom[ 122] = 2'b00;
        w1_rom[ 123] = 2'b00;
        w1_rom[ 124] = 2'b00;
        w1_rom[ 125] = 2'b11;
        w1_rom[ 126] = 2'b01;
        w1_rom[ 127] = 2'b00;
        // Weights  128- 143
        w1_rom[ 128] = 2'b00;
        w1_rom[ 129] = 2'b00;
        w1_rom[ 130] = 2'b01;
        w1_rom[ 131] = 2'b01;
        w1_rom[ 132] = 2'b01;
        w1_rom[ 133] = 2'b00;
        w1_rom[ 134] = 2'b01;
        w1_rom[ 135] = 2'b00;
        w1_rom[ 136] = 2'b00;
        w1_rom[ 137] = 2'b00;
        w1_rom[ 138] = 2'b00;
        w1_rom[ 139] = 2'b00;
        w1_rom[ 140] = 2'b00;
        w1_rom[ 141] = 2'b00;
        w1_rom[ 142] = 2'b11;
        w1_rom[ 143] = 2'b11;
        // Weights  144- 159
        w1_rom[ 144] = 2'b01;
        w1_rom[ 145] = 2'b01;
        w1_rom[ 146] = 2'b00;
        w1_rom[ 147] = 2'b01;
        w1_rom[ 148] = 2'b01;
        w1_rom[ 149] = 2'b00;
        w1_rom[ 150] = 2'b00;
        w1_rom[ 151] = 2'b11;
        w1_rom[ 152] = 2'b01;
        w1_rom[ 153] = 2'b01;
        w1_rom[ 154] = 2'b00;
        w1_rom[ 155] = 2'b11;
        w1_rom[ 156] = 2'b11;
        w1_rom[ 157] = 2'b01;
        w1_rom[ 158] = 2'b01;
        w1_rom[ 159] = 2'b11;
        // Weights  160- 175
        w1_rom[ 160] = 2'b11;
        w1_rom[ 161] = 2'b00;
        w1_rom[ 162] = 2'b00;
        w1_rom[ 163] = 2'b11;
        w1_rom[ 164] = 2'b00;
        w1_rom[ 165] = 2'b00;
        w1_rom[ 166] = 2'b00;
        w1_rom[ 167] = 2'b00;
        w1_rom[ 168] = 2'b00;
        w1_rom[ 169] = 2'b11;
        w1_rom[ 170] = 2'b01;
        w1_rom[ 171] = 2'b01;
        w1_rom[ 172] = 2'b00;
        w1_rom[ 173] = 2'b00;
        w1_rom[ 174] = 2'b00;
        w1_rom[ 175] = 2'b00;
        // Weights  176- 191
        w1_rom[ 176] = 2'b00;
        w1_rom[ 177] = 2'b00;
        w1_rom[ 178] = 2'b00;
        w1_rom[ 179] = 2'b00;
        w1_rom[ 180] = 2'b11;
        w1_rom[ 181] = 2'b11;
        w1_rom[ 182] = 2'b11;
        w1_rom[ 183] = 2'b01;
        w1_rom[ 184] = 2'b00;
        w1_rom[ 185] = 2'b00;
        w1_rom[ 186] = 2'b01;
        w1_rom[ 187] = 2'b01;
        w1_rom[ 188] = 2'b01;
        w1_rom[ 189] = 2'b01;
        w1_rom[ 190] = 2'b01;
        w1_rom[ 191] = 2'b00;
        // Weights  192- 207
        w1_rom[ 192] = 2'b00;
        w1_rom[ 193] = 2'b00;
        w1_rom[ 194] = 2'b00;
        w1_rom[ 195] = 2'b11;
        w1_rom[ 196] = 2'b00;
        w1_rom[ 197] = 2'b01;
        w1_rom[ 198] = 2'b00;
        w1_rom[ 199] = 2'b11;
        w1_rom[ 200] = 2'b00;
        w1_rom[ 201] = 2'b00;
        w1_rom[ 202] = 2'b00;
        w1_rom[ 203] = 2'b11;
        w1_rom[ 204] = 2'b11;
        w1_rom[ 205] = 2'b00;
        w1_rom[ 206] = 2'b01;
        w1_rom[ 207] = 2'b01;
        // Weights  208- 223
        w1_rom[ 208] = 2'b11;
        w1_rom[ 209] = 2'b11;
        w1_rom[ 210] = 2'b11;
        w1_rom[ 211] = 2'b01;
        w1_rom[ 212] = 2'b11;
        w1_rom[ 213] = 2'b11;
        w1_rom[ 214] = 2'b11;
        w1_rom[ 215] = 2'b01;
        w1_rom[ 216] = 2'b11;
        w1_rom[ 217] = 2'b11;
        w1_rom[ 218] = 2'b01;
        w1_rom[ 219] = 2'b00;
        w1_rom[ 220] = 2'b11;
        w1_rom[ 221] = 2'b00;
        w1_rom[ 222] = 2'b11;
        w1_rom[ 223] = 2'b11;
        // Weights  224- 239
        w1_rom[ 224] = 2'b00;
        w1_rom[ 225] = 2'b00;
        w1_rom[ 226] = 2'b01;
        w1_rom[ 227] = 2'b01;
        w1_rom[ 228] = 2'b01;
        w1_rom[ 229] = 2'b01;
        w1_rom[ 230] = 2'b11;
        w1_rom[ 231] = 2'b11;
        w1_rom[ 232] = 2'b11;
        w1_rom[ 233] = 2'b11;
        w1_rom[ 234] = 2'b11;
        w1_rom[ 235] = 2'b11;
        w1_rom[ 236] = 2'b01;
        w1_rom[ 237] = 2'b01;
        w1_rom[ 238] = 2'b00;
        w1_rom[ 239] = 2'b00;
        // Weights  240- 255
        w1_rom[ 240] = 2'b11;
        w1_rom[ 241] = 2'b11;
        w1_rom[ 242] = 2'b11;
        w1_rom[ 243] = 2'b11;
        w1_rom[ 244] = 2'b11;
        w1_rom[ 245] = 2'b01;
        w1_rom[ 246] = 2'b01;
        w1_rom[ 247] = 2'b01;
        w1_rom[ 248] = 2'b00;
        w1_rom[ 249] = 2'b00;
        w1_rom[ 250] = 2'b00;
        w1_rom[ 251] = 2'b11;
        w1_rom[ 252] = 2'b11;
        w1_rom[ 253] = 2'b01;
        w1_rom[ 254] = 2'b01;
        w1_rom[ 255] = 2'b00;

        // Weights  256- 271
        w1_rom[ 256] = 2'b01;
        w1_rom[ 257] = 2'b11;
        w1_rom[ 258] = 2'b11;
        w1_rom[ 259] = 2'b00;
        w1_rom[ 260] = 2'b11;
        w1_rom[ 261] = 2'b00;
        w1_rom[ 262] = 2'b00;
        w1_rom[ 263] = 2'b00;
        w1_rom[ 264] = 2'b11;
        w1_rom[ 265] = 2'b11;
        w1_rom[ 266] = 2'b11;
        w1_rom[ 267] = 2'b11;
        w1_rom[ 268] = 2'b00;
        w1_rom[ 269] = 2'b11;
        w1_rom[ 270] = 2'b00;
        w1_rom[ 271] = 2'b00;
        // Weights  272- 287
        w1_rom[ 272] = 2'b00;
        w1_rom[ 273] = 2'b01;
        w1_rom[ 274] = 2'b00;
        w1_rom[ 275] = 2'b01;
        w1_rom[ 276] = 2'b01;
        w1_rom[ 277] = 2'b01;
        w1_rom[ 278] = 2'b11;
        w1_rom[ 279] = 2'b11;
        w1_rom[ 280] = 2'b01;
        w1_rom[ 281] = 2'b01;
        w1_rom[ 282] = 2'b01;
        w1_rom[ 283] = 2'b11;
        w1_rom[ 284] = 2'b00;
        w1_rom[ 285] = 2'b01;
        w1_rom[ 286] = 2'b01;
        w1_rom[ 287] = 2'b00;
        // Weights  288- 303
        w1_rom[ 288] = 2'b11;
        w1_rom[ 289] = 2'b00;
        w1_rom[ 290] = 2'b11;
        w1_rom[ 291] = 2'b11;
        w1_rom[ 292] = 2'b11;
        w1_rom[ 293] = 2'b11;
        w1_rom[ 294] = 2'b11;
        w1_rom[ 295] = 2'b00;
        w1_rom[ 296] = 2'b00;
        w1_rom[ 297] = 2'b11;
        w1_rom[ 298] = 2'b11;
        w1_rom[ 299] = 2'b01;
        w1_rom[ 300] = 2'b00;
        w1_rom[ 301] = 2'b11;
        w1_rom[ 302] = 2'b11;
        w1_rom[ 303] = 2'b01;
        // Weights  304- 319
        w1_rom[ 304] = 2'b00;
        w1_rom[ 305] = 2'b11;
        w1_rom[ 306] = 2'b00;
        w1_rom[ 307] = 2'b11;
        w1_rom[ 308] = 2'b00;
        w1_rom[ 309] = 2'b11;
        w1_rom[ 310] = 2'b11;
        w1_rom[ 311] = 2'b00;
        w1_rom[ 312] = 2'b11;
        w1_rom[ 313] = 2'b00;
        w1_rom[ 314] = 2'b01;
        w1_rom[ 315] = 2'b00;
        w1_rom[ 316] = 2'b01;
        w1_rom[ 317] = 2'b01;
        w1_rom[ 318] = 2'b01;
        w1_rom[ 319] = 2'b11;
        // Weights  320- 335
        w1_rom[ 320] = 2'b01;
        w1_rom[ 321] = 2'b00;
        w1_rom[ 322] = 2'b11;
        w1_rom[ 323] = 2'b11;
        w1_rom[ 324] = 2'b11;
        w1_rom[ 325] = 2'b11;
        w1_rom[ 326] = 2'b00;
        w1_rom[ 327] = 2'b01;
        w1_rom[ 328] = 2'b00;
        w1_rom[ 329] = 2'b11;
        w1_rom[ 330] = 2'b01;
        w1_rom[ 331] = 2'b00;
        w1_rom[ 332] = 2'b00;
        w1_rom[ 333] = 2'b00;
        w1_rom[ 334] = 2'b01;
        w1_rom[ 335] = 2'b00;
        // Weights  336- 351
        w1_rom[ 336] = 2'b00;
        w1_rom[ 337] = 2'b00;
        w1_rom[ 338] = 2'b01;
        w1_rom[ 339] = 2'b00;
        w1_rom[ 340] = 2'b11;
        w1_rom[ 341] = 2'b00;
        w1_rom[ 342] = 2'b00;
        w1_rom[ 343] = 2'b11;
        w1_rom[ 344] = 2'b00;
        w1_rom[ 345] = 2'b11;
        w1_rom[ 346] = 2'b11;
        w1_rom[ 347] = 2'b11;
        w1_rom[ 348] = 2'b11;
        w1_rom[ 349] = 2'b00;
        w1_rom[ 350] = 2'b11;
        w1_rom[ 351] = 2'b11;
        // Weights  352- 367
        w1_rom[ 352] = 2'b00;
        w1_rom[ 353] = 2'b11;
        w1_rom[ 354] = 2'b01;
        w1_rom[ 355] = 2'b00;
        w1_rom[ 356] = 2'b01;
        w1_rom[ 357] = 2'b00;
        w1_rom[ 358] = 2'b11;
        w1_rom[ 359] = 2'b01;
        w1_rom[ 360] = 2'b00;
        w1_rom[ 361] = 2'b01;
        w1_rom[ 362] = 2'b00;
        w1_rom[ 363] = 2'b01;
        w1_rom[ 364] = 2'b01;
        w1_rom[ 365] = 2'b00;
        w1_rom[ 366] = 2'b01;
        w1_rom[ 367] = 2'b01;
        // Weights  368- 383
        w1_rom[ 368] = 2'b00;
        w1_rom[ 369] = 2'b00;
        w1_rom[ 370] = 2'b00;
        w1_rom[ 371] = 2'b11;
        w1_rom[ 372] = 2'b11;
        w1_rom[ 373] = 2'b01;
        w1_rom[ 374] = 2'b01;
        w1_rom[ 375] = 2'b01;
        w1_rom[ 376] = 2'b00;
        w1_rom[ 377] = 2'b11;
        w1_rom[ 378] = 2'b11;
        w1_rom[ 379] = 2'b11;
        w1_rom[ 380] = 2'b11;
        w1_rom[ 381] = 2'b11;
        w1_rom[ 382] = 2'b00;
        w1_rom[ 383] = 2'b11;
        // Weights  384- 399
        w1_rom[ 384] = 2'b00;
        w1_rom[ 385] = 2'b01;
        w1_rom[ 386] = 2'b00;
        w1_rom[ 387] = 2'b01;
        w1_rom[ 388] = 2'b01;
        w1_rom[ 389] = 2'b01;
        w1_rom[ 390] = 2'b00;
        w1_rom[ 391] = 2'b11;
        w1_rom[ 392] = 2'b00;
        w1_rom[ 393] = 2'b00;
        w1_rom[ 394] = 2'b11;
        w1_rom[ 395] = 2'b11;
        w1_rom[ 396] = 2'b11;
        w1_rom[ 397] = 2'b01;
        w1_rom[ 398] = 2'b01;
        w1_rom[ 399] = 2'b00;
        // Weights  400- 415
        w1_rom[ 400] = 2'b00;
        w1_rom[ 401] = 2'b00;
        w1_rom[ 402] = 2'b01;
        w1_rom[ 403] = 2'b11;
        w1_rom[ 404] = 2'b11;
        w1_rom[ 405] = 2'b11;
        w1_rom[ 406] = 2'b11;
        w1_rom[ 407] = 2'b01;
        w1_rom[ 408] = 2'b00;
        w1_rom[ 409] = 2'b01;
        w1_rom[ 410] = 2'b01;
        w1_rom[ 411] = 2'b01;
        w1_rom[ 412] = 2'b00;
        w1_rom[ 413] = 2'b11;
        w1_rom[ 414] = 2'b01;
        w1_rom[ 415] = 2'b00;
        // Weights  416- 431
        w1_rom[ 416] = 2'b00;
        w1_rom[ 417] = 2'b00;
        w1_rom[ 418] = 2'b00;
        w1_rom[ 419] = 2'b01;
        w1_rom[ 420] = 2'b11;
        w1_rom[ 421] = 2'b11;
        w1_rom[ 422] = 2'b01;
        w1_rom[ 423] = 2'b11;
        w1_rom[ 424] = 2'b11;
        w1_rom[ 425] = 2'b11;
        w1_rom[ 426] = 2'b00;
        w1_rom[ 427] = 2'b01;
        w1_rom[ 428] = 2'b00;
        w1_rom[ 429] = 2'b01;
        w1_rom[ 430] = 2'b00;
        w1_rom[ 431] = 2'b11;
        // Weights  432- 447
        w1_rom[ 432] = 2'b00;
        w1_rom[ 433] = 2'b00;
        w1_rom[ 434] = 2'b00;
        w1_rom[ 435] = 2'b01;
        w1_rom[ 436] = 2'b01;
        w1_rom[ 437] = 2'b00;
        w1_rom[ 438] = 2'b11;
        w1_rom[ 439] = 2'b00;
        w1_rom[ 440] = 2'b00;
        w1_rom[ 441] = 2'b00;
        w1_rom[ 442] = 2'b00;
        w1_rom[ 443] = 2'b11;
        w1_rom[ 444] = 2'b00;
        w1_rom[ 445] = 2'b11;
        w1_rom[ 446] = 2'b11;
        w1_rom[ 447] = 2'b00;
        // Weights  448- 463
        w1_rom[ 448] = 2'b00;
        w1_rom[ 449] = 2'b00;
        w1_rom[ 450] = 2'b00;
        w1_rom[ 451] = 2'b11;
        w1_rom[ 452] = 2'b00;
        w1_rom[ 453] = 2'b11;
        w1_rom[ 454] = 2'b00;
        w1_rom[ 455] = 2'b00;
        w1_rom[ 456] = 2'b00;
        w1_rom[ 457] = 2'b00;
        w1_rom[ 458] = 2'b11;
        w1_rom[ 459] = 2'b00;
        w1_rom[ 460] = 2'b00;
        w1_rom[ 461] = 2'b00;
        w1_rom[ 462] = 2'b00;
        w1_rom[ 463] = 2'b01;
        // Weights  464- 479
        w1_rom[ 464] = 2'b00;
        w1_rom[ 465] = 2'b00;
        w1_rom[ 466] = 2'b00;
        w1_rom[ 467] = 2'b00;
        w1_rom[ 468] = 2'b00;
        w1_rom[ 469] = 2'b01;
        w1_rom[ 470] = 2'b01;
        w1_rom[ 471] = 2'b01;
        w1_rom[ 472] = 2'b00;
        w1_rom[ 473] = 2'b01;
        w1_rom[ 474] = 2'b01;
        w1_rom[ 475] = 2'b01;
        w1_rom[ 476] = 2'b00;
        w1_rom[ 477] = 2'b11;
        w1_rom[ 478] = 2'b11;
        w1_rom[ 479] = 2'b01;
        // Weights  480- 495
        w1_rom[ 480] = 2'b00;
        w1_rom[ 481] = 2'b00;
        w1_rom[ 482] = 2'b00;
        w1_rom[ 483] = 2'b01;
        w1_rom[ 484] = 2'b00;
        w1_rom[ 485] = 2'b00;
        w1_rom[ 486] = 2'b00;
        w1_rom[ 487] = 2'b00;
        w1_rom[ 488] = 2'b00;
        w1_rom[ 489] = 2'b00;
        w1_rom[ 490] = 2'b00;
        w1_rom[ 491] = 2'b11;
        w1_rom[ 492] = 2'b00;
        w1_rom[ 493] = 2'b00;
        w1_rom[ 494] = 2'b00;
        w1_rom[ 495] = 2'b00;
        // Weights  496- 511
        w1_rom[ 496] = 2'b00;
        w1_rom[ 497] = 2'b00;
        w1_rom[ 498] = 2'b00;
        w1_rom[ 499] = 2'b00;
        w1_rom[ 500] = 2'b00;
        w1_rom[ 501] = 2'b00;
        w1_rom[ 502] = 2'b11;
        w1_rom[ 503] = 2'b00;
        w1_rom[ 504] = 2'b00;
        w1_rom[ 505] = 2'b00;
        w1_rom[ 506] = 2'b00;
        w1_rom[ 507] = 2'b00;
        w1_rom[ 508] = 2'b00;
        w1_rom[ 509] = 2'b11;
        w1_rom[ 510] = 2'b00;
        w1_rom[ 511] = 2'b00;

        // Weights  512- 527
        w1_rom[ 512] = 2'b00;
        w1_rom[ 513] = 2'b00;
        w1_rom[ 514] = 2'b11;
        w1_rom[ 515] = 2'b11;
        w1_rom[ 516] = 2'b11;
        w1_rom[ 517] = 2'b11;
        w1_rom[ 518] = 2'b00;
        w1_rom[ 519] = 2'b00;
        w1_rom[ 520] = 2'b00;
        w1_rom[ 521] = 2'b00;
        w1_rom[ 522] = 2'b11;
        w1_rom[ 523] = 2'b11;
        w1_rom[ 524] = 2'b01;
        w1_rom[ 525] = 2'b00;
        w1_rom[ 526] = 2'b01;
        w1_rom[ 527] = 2'b00;
        // Weights  528- 543
        w1_rom[ 528] = 2'b11;
        w1_rom[ 529] = 2'b11;
        w1_rom[ 530] = 2'b01;
        w1_rom[ 531] = 2'b00;
        w1_rom[ 532] = 2'b11;
        w1_rom[ 533] = 2'b00;
        w1_rom[ 534] = 2'b01;
        w1_rom[ 535] = 2'b01;
        w1_rom[ 536] = 2'b00;
        w1_rom[ 537] = 2'b01;
        w1_rom[ 538] = 2'b01;
        w1_rom[ 539] = 2'b01;
        w1_rom[ 540] = 2'b01;
        w1_rom[ 541] = 2'b01;
        w1_rom[ 542] = 2'b11;
        w1_rom[ 543] = 2'b00;
        // Weights  544- 559
        w1_rom[ 544] = 2'b00;
        w1_rom[ 545] = 2'b11;
        w1_rom[ 546] = 2'b11;
        w1_rom[ 547] = 2'b01;
        w1_rom[ 548] = 2'b01;
        w1_rom[ 549] = 2'b00;
        w1_rom[ 550] = 2'b11;
        w1_rom[ 551] = 2'b11;
        w1_rom[ 552] = 2'b00;
        w1_rom[ 553] = 2'b11;
        w1_rom[ 554] = 2'b11;
        w1_rom[ 555] = 2'b11;
        w1_rom[ 556] = 2'b11;
        w1_rom[ 557] = 2'b11;
        w1_rom[ 558] = 2'b11;
        w1_rom[ 559] = 2'b11;
        // Weights  560- 575
        w1_rom[ 560] = 2'b00;
        w1_rom[ 561] = 2'b00;
        w1_rom[ 562] = 2'b00;
        w1_rom[ 563] = 2'b00;
        w1_rom[ 564] = 2'b00;
        w1_rom[ 565] = 2'b01;
        w1_rom[ 566] = 2'b01;
        w1_rom[ 567] = 2'b00;
        w1_rom[ 568] = 2'b01;
        w1_rom[ 569] = 2'b00;
        w1_rom[ 570] = 2'b01;
        w1_rom[ 571] = 2'b01;
        w1_rom[ 572] = 2'b01;
        w1_rom[ 573] = 2'b01;
        w1_rom[ 574] = 2'b01;
        w1_rom[ 575] = 2'b00;
        // Weights  576- 591
        w1_rom[ 576] = 2'b00;
        w1_rom[ 577] = 2'b00;
        w1_rom[ 578] = 2'b00;
        w1_rom[ 579] = 2'b00;
        w1_rom[ 580] = 2'b11;
        w1_rom[ 581] = 2'b11;
        w1_rom[ 582] = 2'b00;
        w1_rom[ 583] = 2'b00;
        w1_rom[ 584] = 2'b00;
        w1_rom[ 585] = 2'b00;
        w1_rom[ 586] = 2'b11;
        w1_rom[ 587] = 2'b11;
        w1_rom[ 588] = 2'b11;
        w1_rom[ 589] = 2'b11;
        w1_rom[ 590] = 2'b11;
        w1_rom[ 591] = 2'b11;
        // Weights  592- 607
        w1_rom[ 592] = 2'b01;
        w1_rom[ 593] = 2'b01;
        w1_rom[ 594] = 2'b00;
        w1_rom[ 595] = 2'b01;
        w1_rom[ 596] = 2'b01;
        w1_rom[ 597] = 2'b01;
        w1_rom[ 598] = 2'b11;
        w1_rom[ 599] = 2'b11;
        w1_rom[ 600] = 2'b01;
        w1_rom[ 601] = 2'b01;
        w1_rom[ 602] = 2'b01;
        w1_rom[ 603] = 2'b11;
        w1_rom[ 604] = 2'b01;
        w1_rom[ 605] = 2'b01;
        w1_rom[ 606] = 2'b01;
        w1_rom[ 607] = 2'b11;
        // Weights  608- 623
        w1_rom[ 608] = 2'b00;
        w1_rom[ 609] = 2'b01;
        w1_rom[ 610] = 2'b11;
        w1_rom[ 611] = 2'b11;
        w1_rom[ 612] = 2'b01;
        w1_rom[ 613] = 2'b01;
        w1_rom[ 614] = 2'b11;
        w1_rom[ 615] = 2'b11;
        w1_rom[ 616] = 2'b00;
        w1_rom[ 617] = 2'b11;
        w1_rom[ 618] = 2'b00;
        w1_rom[ 619] = 2'b11;
        w1_rom[ 620] = 2'b00;
        w1_rom[ 621] = 2'b11;
        w1_rom[ 622] = 2'b11;
        w1_rom[ 623] = 2'b11;
        // Weights  624- 639
        w1_rom[ 624] = 2'b00;
        w1_rom[ 625] = 2'b11;
        w1_rom[ 626] = 2'b11;
        w1_rom[ 627] = 2'b00;
        w1_rom[ 628] = 2'b00;
        w1_rom[ 629] = 2'b11;
        w1_rom[ 630] = 2'b11;
        w1_rom[ 631] = 2'b00;
        w1_rom[ 632] = 2'b00;
        w1_rom[ 633] = 2'b01;
        w1_rom[ 634] = 2'b01;
        w1_rom[ 635] = 2'b01;
        w1_rom[ 636] = 2'b01;
        w1_rom[ 637] = 2'b01;
        w1_rom[ 638] = 2'b01;
        w1_rom[ 639] = 2'b01;
        // Weights  640- 655
        w1_rom[ 640] = 2'b11;
        w1_rom[ 641] = 2'b11;
        w1_rom[ 642] = 2'b00;
        w1_rom[ 643] = 2'b11;
        w1_rom[ 644] = 2'b11;
        w1_rom[ 645] = 2'b00;
        w1_rom[ 646] = 2'b11;
        w1_rom[ 647] = 2'b00;
        w1_rom[ 648] = 2'b00;
        w1_rom[ 649] = 2'b01;
        w1_rom[ 650] = 2'b00;
        w1_rom[ 651] = 2'b00;
        w1_rom[ 652] = 2'b11;
        w1_rom[ 653] = 2'b00;
        w1_rom[ 654] = 2'b01;
        w1_rom[ 655] = 2'b00;
        // Weights  656- 671
        w1_rom[ 656] = 2'b00;
        w1_rom[ 657] = 2'b00;
        w1_rom[ 658] = 2'b00;
        w1_rom[ 659] = 2'b11;
        w1_rom[ 660] = 2'b11;
        w1_rom[ 661] = 2'b01;
        w1_rom[ 662] = 2'b01;
        w1_rom[ 663] = 2'b01;
        w1_rom[ 664] = 2'b00;
        w1_rom[ 665] = 2'b11;
        w1_rom[ 666] = 2'b11;
        w1_rom[ 667] = 2'b01;
        w1_rom[ 668] = 2'b01;
        w1_rom[ 669] = 2'b11;
        w1_rom[ 670] = 2'b11;
        w1_rom[ 671] = 2'b00;
        // Weights  672- 687
        w1_rom[ 672] = 2'b00;
        w1_rom[ 673] = 2'b01;
        w1_rom[ 674] = 2'b01;
        w1_rom[ 675] = 2'b01;
        w1_rom[ 676] = 2'b00;
        w1_rom[ 677] = 2'b01;
        w1_rom[ 678] = 2'b00;
        w1_rom[ 679] = 2'b00;
        w1_rom[ 680] = 2'b00;
        w1_rom[ 681] = 2'b01;
        w1_rom[ 682] = 2'b11;
        w1_rom[ 683] = 2'b11;
        w1_rom[ 684] = 2'b00;
        w1_rom[ 685] = 2'b00;
        w1_rom[ 686] = 2'b00;
        w1_rom[ 687] = 2'b00;
        // Weights  688- 703
        w1_rom[ 688] = 2'b00;
        w1_rom[ 689] = 2'b00;
        w1_rom[ 690] = 2'b00;
        w1_rom[ 691] = 2'b11;
        w1_rom[ 692] = 2'b00;
        w1_rom[ 693] = 2'b01;
        w1_rom[ 694] = 2'b01;
        w1_rom[ 695] = 2'b00;
        w1_rom[ 696] = 2'b00;
        w1_rom[ 697] = 2'b00;
        w1_rom[ 698] = 2'b00;
        w1_rom[ 699] = 2'b11;
        w1_rom[ 700] = 2'b11;
        w1_rom[ 701] = 2'b11;
        w1_rom[ 702] = 2'b00;
        w1_rom[ 703] = 2'b00;
        // Weights  704- 719
        w1_rom[ 704] = 2'b11;
        w1_rom[ 705] = 2'b01;
        w1_rom[ 706] = 2'b11;
        w1_rom[ 707] = 2'b11;
        w1_rom[ 708] = 2'b11;
        w1_rom[ 709] = 2'b00;
        w1_rom[ 710] = 2'b00;
        w1_rom[ 711] = 2'b00;
        w1_rom[ 712] = 2'b00;
        w1_rom[ 713] = 2'b00;
        w1_rom[ 714] = 2'b11;
        w1_rom[ 715] = 2'b11;
        w1_rom[ 716] = 2'b11;
        w1_rom[ 717] = 2'b00;
        w1_rom[ 718] = 2'b01;
        w1_rom[ 719] = 2'b01;
        // Weights  720- 735
        w1_rom[ 720] = 2'b11;
        w1_rom[ 721] = 2'b11;
        w1_rom[ 722] = 2'b01;
        w1_rom[ 723] = 2'b00;
        w1_rom[ 724] = 2'b11;
        w1_rom[ 725] = 2'b00;
        w1_rom[ 726] = 2'b01;
        w1_rom[ 727] = 2'b01;
        w1_rom[ 728] = 2'b00;
        w1_rom[ 729] = 2'b11;
        w1_rom[ 730] = 2'b00;
        w1_rom[ 731] = 2'b01;
        w1_rom[ 732] = 2'b11;
        w1_rom[ 733] = 2'b11;
        w1_rom[ 734] = 2'b11;
        w1_rom[ 735] = 2'b00;
        // Weights  736- 751
        w1_rom[ 736] = 2'b00;
        w1_rom[ 737] = 2'b01;
        w1_rom[ 738] = 2'b00;
        w1_rom[ 739] = 2'b11;
        w1_rom[ 740] = 2'b00;
        w1_rom[ 741] = 2'b01;
        w1_rom[ 742] = 2'b00;
        w1_rom[ 743] = 2'b00;
        w1_rom[ 744] = 2'b00;
        w1_rom[ 745] = 2'b00;
        w1_rom[ 746] = 2'b11;
        w1_rom[ 747] = 2'b11;
        w1_rom[ 748] = 2'b01;
        w1_rom[ 749] = 2'b11;
        w1_rom[ 750] = 2'b11;
        w1_rom[ 751] = 2'b00;
        // Weights  752- 767
        w1_rom[ 752] = 2'b11;
        w1_rom[ 753] = 2'b11;
        w1_rom[ 754] = 2'b00;
        w1_rom[ 755] = 2'b00;
        w1_rom[ 756] = 2'b00;
        w1_rom[ 757] = 2'b01;
        w1_rom[ 758] = 2'b01;
        w1_rom[ 759] = 2'b00;
        w1_rom[ 760] = 2'b00;
        w1_rom[ 761] = 2'b00;
        w1_rom[ 762] = 2'b11;
        w1_rom[ 763] = 2'b11;
        w1_rom[ 764] = 2'b11;
        w1_rom[ 765] = 2'b11;
        w1_rom[ 766] = 2'b00;
        w1_rom[ 767] = 2'b00;

        // Weights  768- 783
        w1_rom[ 768] = 2'b11;
        w1_rom[ 769] = 2'b00;
        w1_rom[ 770] = 2'b00;
        w1_rom[ 771] = 2'b00;
        w1_rom[ 772] = 2'b00;
        w1_rom[ 773] = 2'b00;
        w1_rom[ 774] = 2'b11;
        w1_rom[ 775] = 2'b00;
        w1_rom[ 776] = 2'b00;
        w1_rom[ 777] = 2'b01;
        w1_rom[ 778] = 2'b00;
        w1_rom[ 779] = 2'b01;
        w1_rom[ 780] = 2'b00;
        w1_rom[ 781] = 2'b00;
        w1_rom[ 782] = 2'b01;
        w1_rom[ 783] = 2'b01;
        // Weights  784- 799
        w1_rom[ 784] = 2'b00;
        w1_rom[ 785] = 2'b11;
        w1_rom[ 786] = 2'b11;
        w1_rom[ 787] = 2'b11;
        w1_rom[ 788] = 2'b01;
        w1_rom[ 789] = 2'b11;
        w1_rom[ 790] = 2'b11;
        w1_rom[ 791] = 2'b01;
        w1_rom[ 792] = 2'b11;
        w1_rom[ 793] = 2'b11;
        w1_rom[ 794] = 2'b11;
        w1_rom[ 795] = 2'b11;
        w1_rom[ 796] = 2'b01;
        w1_rom[ 797] = 2'b11;
        w1_rom[ 798] = 2'b11;
        w1_rom[ 799] = 2'b00;
        // Weights  800- 815
        w1_rom[ 800] = 2'b11;
        w1_rom[ 801] = 2'b11;
        w1_rom[ 802] = 2'b11;
        w1_rom[ 803] = 2'b01;
        w1_rom[ 804] = 2'b01;
        w1_rom[ 805] = 2'b00;
        w1_rom[ 806] = 2'b11;
        w1_rom[ 807] = 2'b11;
        w1_rom[ 808] = 2'b00;
        w1_rom[ 809] = 2'b01;
        w1_rom[ 810] = 2'b11;
        w1_rom[ 811] = 2'b11;
        w1_rom[ 812] = 2'b01;
        w1_rom[ 813] = 2'b01;
        w1_rom[ 814] = 2'b01;
        w1_rom[ 815] = 2'b00;
        // Weights  816- 831
        w1_rom[ 816] = 2'b00;
        w1_rom[ 817] = 2'b01;
        w1_rom[ 818] = 2'b01;
        w1_rom[ 819] = 2'b11;
        w1_rom[ 820] = 2'b00;
        w1_rom[ 821] = 2'b01;
        w1_rom[ 822] = 2'b01;
        w1_rom[ 823] = 2'b00;
        w1_rom[ 824] = 2'b00;
        w1_rom[ 825] = 2'b00;
        w1_rom[ 826] = 2'b00;
        w1_rom[ 827] = 2'b11;
        w1_rom[ 828] = 2'b11;
        w1_rom[ 829] = 2'b11;
        w1_rom[ 830] = 2'b00;
        w1_rom[ 831] = 2'b00;
        // Weights  832- 847
        w1_rom[ 832] = 2'b00;
        w1_rom[ 833] = 2'b00;
        w1_rom[ 834] = 2'b00;
        w1_rom[ 835] = 2'b11;
        w1_rom[ 836] = 2'b01;
        w1_rom[ 837] = 2'b00;
        w1_rom[ 838] = 2'b11;
        w1_rom[ 839] = 2'b00;
        w1_rom[ 840] = 2'b11;
        w1_rom[ 841] = 2'b00;
        w1_rom[ 842] = 2'b00;
        w1_rom[ 843] = 2'b11;
        w1_rom[ 844] = 2'b11;
        w1_rom[ 845] = 2'b00;
        w1_rom[ 846] = 2'b00;
        w1_rom[ 847] = 2'b00;
        // Weights  848- 863
        w1_rom[ 848] = 2'b00;
        w1_rom[ 849] = 2'b01;
        w1_rom[ 850] = 2'b00;
        w1_rom[ 851] = 2'b11;
        w1_rom[ 852] = 2'b11;
        w1_rom[ 853] = 2'b00;
        w1_rom[ 854] = 2'b01;
        w1_rom[ 855] = 2'b11;
        w1_rom[ 856] = 2'b01;
        w1_rom[ 857] = 2'b00;
        w1_rom[ 858] = 2'b11;
        w1_rom[ 859] = 2'b00;
        w1_rom[ 860] = 2'b01;
        w1_rom[ 861] = 2'b01;
        w1_rom[ 862] = 2'b01;
        w1_rom[ 863] = 2'b00;
        // Weights  864- 879
        w1_rom[ 864] = 2'b00;
        w1_rom[ 865] = 2'b01;
        w1_rom[ 866] = 2'b00;
        w1_rom[ 867] = 2'b11;
        w1_rom[ 868] = 2'b00;
        w1_rom[ 869] = 2'b01;
        w1_rom[ 870] = 2'b01;
        w1_rom[ 871] = 2'b01;
        w1_rom[ 872] = 2'b00;
        w1_rom[ 873] = 2'b11;
        w1_rom[ 874] = 2'b00;
        w1_rom[ 875] = 2'b01;
        w1_rom[ 876] = 2'b00;
        w1_rom[ 877] = 2'b00;
        w1_rom[ 878] = 2'b11;
        w1_rom[ 879] = 2'b00;
        // Weights  880- 895
        w1_rom[ 880] = 2'b00;
        w1_rom[ 881] = 2'b00;
        w1_rom[ 882] = 2'b11;
        w1_rom[ 883] = 2'b00;
        w1_rom[ 884] = 2'b01;
        w1_rom[ 885] = 2'b01;
        w1_rom[ 886] = 2'b11;
        w1_rom[ 887] = 2'b01;
        w1_rom[ 888] = 2'b11;
        w1_rom[ 889] = 2'b01;
        w1_rom[ 890] = 2'b11;
        w1_rom[ 891] = 2'b11;
        w1_rom[ 892] = 2'b00;
        w1_rom[ 893] = 2'b11;
        w1_rom[ 894] = 2'b11;
        w1_rom[ 895] = 2'b00;
        // Weights  896- 911
        w1_rom[ 896] = 2'b00;
        w1_rom[ 897] = 2'b00;
        w1_rom[ 898] = 2'b00;
        w1_rom[ 899] = 2'b00;
        w1_rom[ 900] = 2'b01;
        w1_rom[ 901] = 2'b01;
        w1_rom[ 902] = 2'b00;
        w1_rom[ 903] = 2'b00;
        w1_rom[ 904] = 2'b00;
        w1_rom[ 905] = 2'b01;
        w1_rom[ 906] = 2'b01;
        w1_rom[ 907] = 2'b00;
        w1_rom[ 908] = 2'b00;
        w1_rom[ 909] = 2'b01;
        w1_rom[ 910] = 2'b01;
        w1_rom[ 911] = 2'b01;
        // Weights  912- 927
        w1_rom[ 912] = 2'b00;
        w1_rom[ 913] = 2'b01;
        w1_rom[ 914] = 2'b11;
        w1_rom[ 915] = 2'b11;
        w1_rom[ 916] = 2'b00;
        w1_rom[ 917] = 2'b11;
        w1_rom[ 918] = 2'b11;
        w1_rom[ 919] = 2'b00;
        w1_rom[ 920] = 2'b00;
        w1_rom[ 921] = 2'b01;
        w1_rom[ 922] = 2'b00;
        w1_rom[ 923] = 2'b01;
        w1_rom[ 924] = 2'b01;
        w1_rom[ 925] = 2'b01;
        w1_rom[ 926] = 2'b11;
        w1_rom[ 927] = 2'b11;
        // Weights  928- 943
        w1_rom[ 928] = 2'b00;
        w1_rom[ 929] = 2'b00;
        w1_rom[ 930] = 2'b00;
        w1_rom[ 931] = 2'b00;
        w1_rom[ 932] = 2'b01;
        w1_rom[ 933] = 2'b01;
        w1_rom[ 934] = 2'b01;
        w1_rom[ 935] = 2'b11;
        w1_rom[ 936] = 2'b00;
        w1_rom[ 937] = 2'b11;
        w1_rom[ 938] = 2'b11;
        w1_rom[ 939] = 2'b11;
        w1_rom[ 940] = 2'b11;
        w1_rom[ 941] = 2'b00;
        w1_rom[ 942] = 2'b11;
        w1_rom[ 943] = 2'b11;
        // Weights  944- 959
        w1_rom[ 944] = 2'b00;
        w1_rom[ 945] = 2'b00;
        w1_rom[ 946] = 2'b00;
        w1_rom[ 947] = 2'b11;
        w1_rom[ 948] = 2'b01;
        w1_rom[ 949] = 2'b00;
        w1_rom[ 950] = 2'b11;
        w1_rom[ 951] = 2'b00;
        w1_rom[ 952] = 2'b00;
        w1_rom[ 953] = 2'b01;
        w1_rom[ 954] = 2'b01;
        w1_rom[ 955] = 2'b01;
        w1_rom[ 956] = 2'b11;
        w1_rom[ 957] = 2'b00;
        w1_rom[ 958] = 2'b00;
        w1_rom[ 959] = 2'b11;
        // Weights  960- 975
        w1_rom[ 960] = 2'b01;
        w1_rom[ 961] = 2'b00;
        w1_rom[ 962] = 2'b00;
        w1_rom[ 963] = 2'b00;
        w1_rom[ 964] = 2'b00;
        w1_rom[ 965] = 2'b01;
        w1_rom[ 966] = 2'b00;
        w1_rom[ 967] = 2'b00;
        w1_rom[ 968] = 2'b00;
        w1_rom[ 969] = 2'b00;
        w1_rom[ 970] = 2'b01;
        w1_rom[ 971] = 2'b11;
        w1_rom[ 972] = 2'b11;
        w1_rom[ 973] = 2'b11;
        w1_rom[ 974] = 2'b11;
        w1_rom[ 975] = 2'b00;
        // Weights  976- 991
        w1_rom[ 976] = 2'b01;
        w1_rom[ 977] = 2'b01;
        w1_rom[ 978] = 2'b01;
        w1_rom[ 979] = 2'b01;
        w1_rom[ 980] = 2'b11;
        w1_rom[ 981] = 2'b11;
        w1_rom[ 982] = 2'b11;
        w1_rom[ 983] = 2'b11;
        w1_rom[ 984] = 2'b01;
        w1_rom[ 985] = 2'b01;
        w1_rom[ 986] = 2'b01;
        w1_rom[ 987] = 2'b11;
        w1_rom[ 988] = 2'b11;
        w1_rom[ 989] = 2'b01;
        w1_rom[ 990] = 2'b11;
        w1_rom[ 991] = 2'b11;
        // Weights  992-1007
        w1_rom[ 992] = 2'b00;
        w1_rom[ 993] = 2'b01;
        w1_rom[ 994] = 2'b01;
        w1_rom[ 995] = 2'b11;
        w1_rom[ 996] = 2'b01;
        w1_rom[ 997] = 2'b01;
        w1_rom[ 998] = 2'b01;
        w1_rom[ 999] = 2'b11;
        w1_rom[1000] = 2'b00;
        w1_rom[1001] = 2'b11;
        w1_rom[1002] = 2'b00;
        w1_rom[1003] = 2'b01;
        w1_rom[1004] = 2'b01;
        w1_rom[1005] = 2'b11;
        w1_rom[1006] = 2'b11;
        w1_rom[1007] = 2'b00;
        // Weights 1008-1023
        w1_rom[1008] = 2'b11;
        w1_rom[1009] = 2'b11;
        w1_rom[1010] = 2'b11;
        w1_rom[1011] = 2'b11;
        w1_rom[1012] = 2'b11;
        w1_rom[1013] = 2'b11;
        w1_rom[1014] = 2'b01;
        w1_rom[1015] = 2'b00;
        w1_rom[1016] = 2'b00;
        w1_rom[1017] = 2'b01;
        w1_rom[1018] = 2'b01;
        w1_rom[1019] = 2'b11;
        w1_rom[1020] = 2'b00;
        w1_rom[1021] = 2'b11;
        w1_rom[1022] = 2'b00;
        w1_rom[1023] = 2'b00;

        // Weights 1024-1039
        w1_rom[1024] = 2'b01;
        w1_rom[1025] = 2'b00;
        w1_rom[1026] = 2'b01;
        w1_rom[1027] = 2'b11;
        w1_rom[1028] = 2'b11;
        w1_rom[1029] = 2'b11;
        w1_rom[1030] = 2'b11;
        w1_rom[1031] = 2'b00;
        w1_rom[1032] = 2'b11;
        w1_rom[1033] = 2'b00;
        w1_rom[1034] = 2'b00;
        w1_rom[1035] = 2'b11;
        w1_rom[1036] = 2'b00;
        w1_rom[1037] = 2'b00;
        w1_rom[1038] = 2'b01;
        w1_rom[1039] = 2'b01;
        // Weights 1040-1055
        w1_rom[1040] = 2'b11;
        w1_rom[1041] = 2'b11;
        w1_rom[1042] = 2'b00;
        w1_rom[1043] = 2'b00;
        w1_rom[1044] = 2'b00;
        w1_rom[1045] = 2'b01;
        w1_rom[1046] = 2'b01;
        w1_rom[1047] = 2'b01;
        w1_rom[1048] = 2'b11;
        w1_rom[1049] = 2'b00;
        w1_rom[1050] = 2'b01;
        w1_rom[1051] = 2'b01;
        w1_rom[1052] = 2'b11;
        w1_rom[1053] = 2'b11;
        w1_rom[1054] = 2'b11;
        w1_rom[1055] = 2'b01;
        // Weights 1056-1071
        w1_rom[1056] = 2'b01;
        w1_rom[1057] = 2'b01;
        w1_rom[1058] = 2'b01;
        w1_rom[1059] = 2'b00;
        w1_rom[1060] = 2'b11;
        w1_rom[1061] = 2'b00;
        w1_rom[1062] = 2'b00;
        w1_rom[1063] = 2'b00;
        w1_rom[1064] = 2'b01;
        w1_rom[1065] = 2'b01;
        w1_rom[1066] = 2'b00;
        w1_rom[1067] = 2'b11;
        w1_rom[1068] = 2'b00;
        w1_rom[1069] = 2'b11;
        w1_rom[1070] = 2'b00;
        w1_rom[1071] = 2'b00;
        // Weights 1072-1087
        w1_rom[1072] = 2'b11;
        w1_rom[1073] = 2'b00;
        w1_rom[1074] = 2'b01;
        w1_rom[1075] = 2'b00;
        w1_rom[1076] = 2'b11;
        w1_rom[1077] = 2'b01;
        w1_rom[1078] = 2'b01;
        w1_rom[1079] = 2'b00;
        w1_rom[1080] = 2'b01;
        w1_rom[1081] = 2'b00;
        w1_rom[1082] = 2'b11;
        w1_rom[1083] = 2'b11;
        w1_rom[1084] = 2'b11;
        w1_rom[1085] = 2'b11;
        w1_rom[1086] = 2'b11;
        w1_rom[1087] = 2'b00;
        // Weights 1088-1103
        w1_rom[1088] = 2'b00;
        w1_rom[1089] = 2'b00;
        w1_rom[1090] = 2'b00;
        w1_rom[1091] = 2'b11;
        w1_rom[1092] = 2'b11;
        w1_rom[1093] = 2'b11;
        w1_rom[1094] = 2'b11;
        w1_rom[1095] = 2'b00;
        w1_rom[1096] = 2'b00;
        w1_rom[1097] = 2'b01;
        w1_rom[1098] = 2'b00;
        w1_rom[1099] = 2'b01;
        w1_rom[1100] = 2'b11;
        w1_rom[1101] = 2'b00;
        w1_rom[1102] = 2'b11;
        w1_rom[1103] = 2'b00;
        // Weights 1104-1119
        w1_rom[1104] = 2'b00;
        w1_rom[1105] = 2'b01;
        w1_rom[1106] = 2'b11;
        w1_rom[1107] = 2'b00;
        w1_rom[1108] = 2'b01;
        w1_rom[1109] = 2'b00;
        w1_rom[1110] = 2'b00;
        w1_rom[1111] = 2'b01;
        w1_rom[1112] = 2'b01;
        w1_rom[1113] = 2'b01;
        w1_rom[1114] = 2'b11;
        w1_rom[1115] = 2'b11;
        w1_rom[1116] = 2'b01;
        w1_rom[1117] = 2'b11;
        w1_rom[1118] = 2'b11;
        w1_rom[1119] = 2'b01;
        // Weights 1120-1135
        w1_rom[1120] = 2'b01;
        w1_rom[1121] = 2'b11;
        w1_rom[1122] = 2'b11;
        w1_rom[1123] = 2'b11;
        w1_rom[1124] = 2'b11;
        w1_rom[1125] = 2'b00;
        w1_rom[1126] = 2'b00;
        w1_rom[1127] = 2'b00;
        w1_rom[1128] = 2'b00;
        w1_rom[1129] = 2'b01;
        w1_rom[1130] = 2'b11;
        w1_rom[1131] = 2'b11;
        w1_rom[1132] = 2'b00;
        w1_rom[1133] = 2'b01;
        w1_rom[1134] = 2'b01;
        w1_rom[1135] = 2'b01;
        // Weights 1136-1151
        w1_rom[1136] = 2'b00;
        w1_rom[1137] = 2'b01;
        w1_rom[1138] = 2'b01;
        w1_rom[1139] = 2'b00;
        w1_rom[1140] = 2'b00;
        w1_rom[1141] = 2'b01;
        w1_rom[1142] = 2'b11;
        w1_rom[1143] = 2'b00;
        w1_rom[1144] = 2'b00;
        w1_rom[1145] = 2'b00;
        w1_rom[1146] = 2'b01;
        w1_rom[1147] = 2'b01;
        w1_rom[1148] = 2'b00;
        w1_rom[1149] = 2'b00;
        w1_rom[1150] = 2'b00;
        w1_rom[1151] = 2'b00;
        // Weights 1152-1167
        w1_rom[1152] = 2'b00;
        w1_rom[1153] = 2'b00;
        w1_rom[1154] = 2'b00;
        w1_rom[1155] = 2'b00;
        w1_rom[1156] = 2'b00;
        w1_rom[1157] = 2'b00;
        w1_rom[1158] = 2'b00;
        w1_rom[1159] = 2'b00;
        w1_rom[1160] = 2'b00;
        w1_rom[1161] = 2'b00;
        w1_rom[1162] = 2'b00;
        w1_rom[1163] = 2'b01;
        w1_rom[1164] = 2'b01;
        w1_rom[1165] = 2'b00;
        w1_rom[1166] = 2'b11;
        w1_rom[1167] = 2'b00;
        // Weights 1168-1183
        w1_rom[1168] = 2'b11;
        w1_rom[1169] = 2'b11;
        w1_rom[1170] = 2'b01;
        w1_rom[1171] = 2'b01;
        w1_rom[1172] = 2'b01;
        w1_rom[1173] = 2'b11;
        w1_rom[1174] = 2'b00;
        w1_rom[1175] = 2'b00;
        w1_rom[1176] = 2'b00;
        w1_rom[1177] = 2'b00;
        w1_rom[1178] = 2'b00;
        w1_rom[1179] = 2'b11;
        w1_rom[1180] = 2'b11;
        w1_rom[1181] = 2'b01;
        w1_rom[1182] = 2'b01;
        w1_rom[1183] = 2'b01;
        // Weights 1184-1199
        w1_rom[1184] = 2'b11;
        w1_rom[1185] = 2'b11;
        w1_rom[1186] = 2'b11;
        w1_rom[1187] = 2'b01;
        w1_rom[1188] = 2'b01;
        w1_rom[1189] = 2'b11;
        w1_rom[1190] = 2'b11;
        w1_rom[1191] = 2'b00;
        w1_rom[1192] = 2'b00;
        w1_rom[1193] = 2'b01;
        w1_rom[1194] = 2'b01;
        w1_rom[1195] = 2'b01;
        w1_rom[1196] = 2'b00;
        w1_rom[1197] = 2'b11;
        w1_rom[1198] = 2'b01;
        w1_rom[1199] = 2'b01;
        // Weights 1200-1215
        w1_rom[1200] = 2'b11;
        w1_rom[1201] = 2'b11;
        w1_rom[1202] = 2'b00;
        w1_rom[1203] = 2'b11;
        w1_rom[1204] = 2'b00;
        w1_rom[1205] = 2'b00;
        w1_rom[1206] = 2'b01;
        w1_rom[1207] = 2'b01;
        w1_rom[1208] = 2'b00;
        w1_rom[1209] = 2'b11;
        w1_rom[1210] = 2'b11;
        w1_rom[1211] = 2'b01;
        w1_rom[1212] = 2'b01;
        w1_rom[1213] = 2'b01;
        w1_rom[1214] = 2'b01;
        w1_rom[1215] = 2'b00;
        // Weights 1216-1231
        w1_rom[1216] = 2'b01;
        w1_rom[1217] = 2'b00;
        w1_rom[1218] = 2'b11;
        w1_rom[1219] = 2'b11;
        w1_rom[1220] = 2'b11;
        w1_rom[1221] = 2'b11;
        w1_rom[1222] = 2'b00;
        w1_rom[1223] = 2'b11;
        w1_rom[1224] = 2'b00;
        w1_rom[1225] = 2'b00;
        w1_rom[1226] = 2'b00;
        w1_rom[1227] = 2'b01;
        w1_rom[1228] = 2'b00;
        w1_rom[1229] = 2'b00;
        w1_rom[1230] = 2'b00;
        w1_rom[1231] = 2'b00;
        // Weights 1232-1247
        w1_rom[1232] = 2'b00;
        w1_rom[1233] = 2'b00;
        w1_rom[1234] = 2'b11;
        w1_rom[1235] = 2'b01;
        w1_rom[1236] = 2'b01;
        w1_rom[1237] = 2'b01;
        w1_rom[1238] = 2'b00;
        w1_rom[1239] = 2'b01;
        w1_rom[1240] = 2'b00;
        w1_rom[1241] = 2'b00;
        w1_rom[1242] = 2'b00;
        w1_rom[1243] = 2'b11;
        w1_rom[1244] = 2'b01;
        w1_rom[1245] = 2'b11;
        w1_rom[1246] = 2'b11;
        w1_rom[1247] = 2'b11;
        // Weights 1248-1263
        w1_rom[1248] = 2'b00;
        w1_rom[1249] = 2'b00;
        w1_rom[1250] = 2'b00;
        w1_rom[1251] = 2'b11;
        w1_rom[1252] = 2'b11;
        w1_rom[1253] = 2'b01;
        w1_rom[1254] = 2'b11;
        w1_rom[1255] = 2'b00;
        w1_rom[1256] = 2'b00;
        w1_rom[1257] = 2'b01;
        w1_rom[1258] = 2'b11;
        w1_rom[1259] = 2'b11;
        w1_rom[1260] = 2'b00;
        w1_rom[1261] = 2'b11;
        w1_rom[1262] = 2'b01;
        w1_rom[1263] = 2'b01;
        // Weights 1264-1279
        w1_rom[1264] = 2'b00;
        w1_rom[1265] = 2'b00;
        w1_rom[1266] = 2'b01;
        w1_rom[1267] = 2'b11;
        w1_rom[1268] = 2'b00;
        w1_rom[1269] = 2'b00;
        w1_rom[1270] = 2'b01;
        w1_rom[1271] = 2'b00;
        w1_rom[1272] = 2'b01;
        w1_rom[1273] = 2'b00;
        w1_rom[1274] = 2'b01;
        w1_rom[1275] = 2'b00;
        w1_rom[1276] = 2'b11;
        w1_rom[1277] = 2'b00;
        w1_rom[1278] = 2'b00;
        w1_rom[1279] = 2'b11;

        // Weights 1280-1295
        w1_rom[1280] = 2'b00;
        w1_rom[1281] = 2'b00;
        w1_rom[1282] = 2'b01;
        w1_rom[1283] = 2'b01;
        w1_rom[1284] = 2'b01;
        w1_rom[1285] = 2'b01;
        w1_rom[1286] = 2'b00;
        w1_rom[1287] = 2'b11;
        w1_rom[1288] = 2'b00;
        w1_rom[1289] = 2'b11;
        w1_rom[1290] = 2'b11;
        w1_rom[1291] = 2'b00;
        w1_rom[1292] = 2'b01;
        w1_rom[1293] = 2'b01;
        w1_rom[1294] = 2'b01;
        w1_rom[1295] = 2'b00;
        // Weights 1296-1311
        w1_rom[1296] = 2'b11;
        w1_rom[1297] = 2'b11;
        w1_rom[1298] = 2'b11;
        w1_rom[1299] = 2'b11;
        w1_rom[1300] = 2'b11;
        w1_rom[1301] = 2'b11;
        w1_rom[1302] = 2'b11;
        w1_rom[1303] = 2'b11;
        w1_rom[1304] = 2'b11;
        w1_rom[1305] = 2'b11;
        w1_rom[1306] = 2'b00;
        w1_rom[1307] = 2'b11;
        w1_rom[1308] = 2'b11;
        w1_rom[1309] = 2'b11;
        w1_rom[1310] = 2'b11;
        w1_rom[1311] = 2'b11;
        // Weights 1312-1327
        w1_rom[1312] = 2'b00;
        w1_rom[1313] = 2'b01;
        w1_rom[1314] = 2'b01;
        w1_rom[1315] = 2'b01;
        w1_rom[1316] = 2'b01;
        w1_rom[1317] = 2'b11;
        w1_rom[1318] = 2'b00;
        w1_rom[1319] = 2'b01;
        w1_rom[1320] = 2'b11;
        w1_rom[1321] = 2'b11;
        w1_rom[1322] = 2'b01;
        w1_rom[1323] = 2'b01;
        w1_rom[1324] = 2'b01;
        w1_rom[1325] = 2'b01;
        w1_rom[1326] = 2'b01;
        w1_rom[1327] = 2'b01;
        // Weights 1328-1343
        w1_rom[1328] = 2'b01;
        w1_rom[1329] = 2'b11;
        w1_rom[1330] = 2'b01;
        w1_rom[1331] = 2'b11;
        w1_rom[1332] = 2'b00;
        w1_rom[1333] = 2'b01;
        w1_rom[1334] = 2'b01;
        w1_rom[1335] = 2'b00;
        w1_rom[1336] = 2'b01;
        w1_rom[1337] = 2'b11;
        w1_rom[1338] = 2'b11;
        w1_rom[1339] = 2'b11;
        w1_rom[1340] = 2'b11;
        w1_rom[1341] = 2'b11;
        w1_rom[1342] = 2'b00;
        w1_rom[1343] = 2'b01;
        // Weights 1344-1359
        w1_rom[1344] = 2'b00;
        w1_rom[1345] = 2'b01;
        w1_rom[1346] = 2'b01;
        w1_rom[1347] = 2'b11;
        w1_rom[1348] = 2'b00;
        w1_rom[1349] = 2'b00;
        w1_rom[1350] = 2'b00;
        w1_rom[1351] = 2'b00;
        w1_rom[1352] = 2'b00;
        w1_rom[1353] = 2'b00;
        w1_rom[1354] = 2'b11;
        w1_rom[1355] = 2'b00;
        w1_rom[1356] = 2'b00;
        w1_rom[1357] = 2'b11;
        w1_rom[1358] = 2'b00;
        w1_rom[1359] = 2'b11;
        // Weights 1360-1375
        w1_rom[1360] = 2'b00;
        w1_rom[1361] = 2'b00;
        w1_rom[1362] = 2'b00;
        w1_rom[1363] = 2'b00;
        w1_rom[1364] = 2'b01;
        w1_rom[1365] = 2'b01;
        w1_rom[1366] = 2'b11;
        w1_rom[1367] = 2'b11;
        w1_rom[1368] = 2'b00;
        w1_rom[1369] = 2'b11;
        w1_rom[1370] = 2'b11;
        w1_rom[1371] = 2'b11;
        w1_rom[1372] = 2'b11;
        w1_rom[1373] = 2'b11;
        w1_rom[1374] = 2'b01;
        w1_rom[1375] = 2'b00;
        // Weights 1376-1391
        w1_rom[1376] = 2'b00;
        w1_rom[1377] = 2'b01;
        w1_rom[1378] = 2'b01;
        w1_rom[1379] = 2'b11;
        w1_rom[1380] = 2'b11;
        w1_rom[1381] = 2'b11;
        w1_rom[1382] = 2'b00;
        w1_rom[1383] = 2'b01;
        w1_rom[1384] = 2'b00;
        w1_rom[1385] = 2'b01;
        w1_rom[1386] = 2'b00;
        w1_rom[1387] = 2'b01;
        w1_rom[1388] = 2'b01;
        w1_rom[1389] = 2'b11;
        w1_rom[1390] = 2'b01;
        w1_rom[1391] = 2'b01;
        // Weights 1392-1407
        w1_rom[1392] = 2'b00;
        w1_rom[1393] = 2'b00;
        w1_rom[1394] = 2'b01;
        w1_rom[1395] = 2'b00;
        w1_rom[1396] = 2'b00;
        w1_rom[1397] = 2'b01;
        w1_rom[1398] = 2'b01;
        w1_rom[1399] = 2'b01;
        w1_rom[1400] = 2'b00;
        w1_rom[1401] = 2'b11;
        w1_rom[1402] = 2'b11;
        w1_rom[1403] = 2'b11;
        w1_rom[1404] = 2'b11;
        w1_rom[1405] = 2'b00;
        w1_rom[1406] = 2'b11;
        w1_rom[1407] = 2'b00;
        // Weights 1408-1423
        w1_rom[1408] = 2'b00;
        w1_rom[1409] = 2'b00;
        w1_rom[1410] = 2'b00;
        w1_rom[1411] = 2'b00;
        w1_rom[1412] = 2'b11;
        w1_rom[1413] = 2'b00;
        w1_rom[1414] = 2'b00;
        w1_rom[1415] = 2'b00;
        w1_rom[1416] = 2'b01;
        w1_rom[1417] = 2'b01;
        w1_rom[1418] = 2'b00;
        w1_rom[1419] = 2'b00;
        w1_rom[1420] = 2'b00;
        w1_rom[1421] = 2'b00;
        w1_rom[1422] = 2'b11;
        w1_rom[1423] = 2'b00;
        // Weights 1424-1439
        w1_rom[1424] = 2'b00;
        w1_rom[1425] = 2'b00;
        w1_rom[1426] = 2'b00;
        w1_rom[1427] = 2'b11;
        w1_rom[1428] = 2'b00;
        w1_rom[1429] = 2'b00;
        w1_rom[1430] = 2'b11;
        w1_rom[1431] = 2'b11;
        w1_rom[1432] = 2'b00;
        w1_rom[1433] = 2'b00;
        w1_rom[1434] = 2'b00;
        w1_rom[1435] = 2'b01;
        w1_rom[1436] = 2'b01;
        w1_rom[1437] = 2'b00;
        w1_rom[1438] = 2'b01;
        w1_rom[1439] = 2'b00;
        // Weights 1440-1455
        w1_rom[1440] = 2'b00;
        w1_rom[1441] = 2'b01;
        w1_rom[1442] = 2'b01;
        w1_rom[1443] = 2'b01;
        w1_rom[1444] = 2'b11;
        w1_rom[1445] = 2'b00;
        w1_rom[1446] = 2'b01;
        w1_rom[1447] = 2'b11;
        w1_rom[1448] = 2'b00;
        w1_rom[1449] = 2'b00;
        w1_rom[1450] = 2'b11;
        w1_rom[1451] = 2'b11;
        w1_rom[1452] = 2'b00;
        w1_rom[1453] = 2'b00;
        w1_rom[1454] = 2'b11;
        w1_rom[1455] = 2'b11;
        // Weights 1456-1471
        w1_rom[1456] = 2'b01;
        w1_rom[1457] = 2'b00;
        w1_rom[1458] = 2'b00;
        w1_rom[1459] = 2'b01;
        w1_rom[1460] = 2'b01;
        w1_rom[1461] = 2'b00;
        w1_rom[1462] = 2'b11;
        w1_rom[1463] = 2'b00;
        w1_rom[1464] = 2'b00;
        w1_rom[1465] = 2'b00;
        w1_rom[1466] = 2'b00;
        w1_rom[1467] = 2'b11;
        w1_rom[1468] = 2'b11;
        w1_rom[1469] = 2'b11;
        w1_rom[1470] = 2'b11;
        w1_rom[1471] = 2'b00;
        // Weights 1472-1487
        w1_rom[1472] = 2'b00;
        w1_rom[1473] = 2'b00;
        w1_rom[1474] = 2'b00;
        w1_rom[1475] = 2'b01;
        w1_rom[1476] = 2'b01;
        w1_rom[1477] = 2'b01;
        w1_rom[1478] = 2'b00;
        w1_rom[1479] = 2'b01;
        w1_rom[1480] = 2'b00;
        w1_rom[1481] = 2'b11;
        w1_rom[1482] = 2'b11;
        w1_rom[1483] = 2'b00;
        w1_rom[1484] = 2'b01;
        w1_rom[1485] = 2'b00;
        w1_rom[1486] = 2'b00;
        w1_rom[1487] = 2'b00;
        // Weights 1488-1503
        w1_rom[1488] = 2'b00;
        w1_rom[1489] = 2'b11;
        w1_rom[1490] = 2'b00;
        w1_rom[1491] = 2'b01;
        w1_rom[1492] = 2'b00;
        w1_rom[1493] = 2'b11;
        w1_rom[1494] = 2'b00;
        w1_rom[1495] = 2'b01;
        w1_rom[1496] = 2'b00;
        w1_rom[1497] = 2'b01;
        w1_rom[1498] = 2'b01;
        w1_rom[1499] = 2'b01;
        w1_rom[1500] = 2'b11;
        w1_rom[1501] = 2'b11;
        w1_rom[1502] = 2'b01;
        w1_rom[1503] = 2'b01;
        // Weights 1504-1519
        w1_rom[1504] = 2'b11;
        w1_rom[1505] = 2'b11;
        w1_rom[1506] = 2'b00;
        w1_rom[1507] = 2'b01;
        w1_rom[1508] = 2'b11;
        w1_rom[1509] = 2'b11;
        w1_rom[1510] = 2'b11;
        w1_rom[1511] = 2'b01;
        w1_rom[1512] = 2'b00;
        w1_rom[1513] = 2'b00;
        w1_rom[1514] = 2'b01;
        w1_rom[1515] = 2'b01;
        w1_rom[1516] = 2'b00;
        w1_rom[1517] = 2'b00;
        w1_rom[1518] = 2'b00;
        w1_rom[1519] = 2'b01;
        // Weights 1520-1535
        w1_rom[1520] = 2'b01;
        w1_rom[1521] = 2'b11;
        w1_rom[1522] = 2'b00;
        w1_rom[1523] = 2'b01;
        w1_rom[1524] = 2'b00;
        w1_rom[1525] = 2'b00;
        w1_rom[1526] = 2'b01;
        w1_rom[1527] = 2'b01;
        w1_rom[1528] = 2'b00;
        w1_rom[1529] = 2'b11;
        w1_rom[1530] = 2'b11;
        w1_rom[1531] = 2'b00;
        w1_rom[1532] = 2'b01;
        w1_rom[1533] = 2'b01;
        w1_rom[1534] = 2'b00;
        w1_rom[1535] = 2'b00;

        // Weights 1536-1551
        w1_rom[1536] = 2'b01;
        w1_rom[1537] = 2'b01;
        w1_rom[1538] = 2'b11;
        w1_rom[1539] = 2'b11;
        w1_rom[1540] = 2'b11;
        w1_rom[1541] = 2'b11;
        w1_rom[1542] = 2'b00;
        w1_rom[1543] = 2'b00;
        w1_rom[1544] = 2'b00;
        w1_rom[1545] = 2'b01;
        w1_rom[1546] = 2'b01;
        w1_rom[1547] = 2'b01;
        w1_rom[1548] = 2'b01;
        w1_rom[1549] = 2'b01;
        w1_rom[1550] = 2'b11;
        w1_rom[1551] = 2'b01;
        // Weights 1552-1567
        w1_rom[1552] = 2'b00;
        w1_rom[1553] = 2'b01;
        w1_rom[1554] = 2'b01;
        w1_rom[1555] = 2'b01;
        w1_rom[1556] = 2'b01;
        w1_rom[1557] = 2'b01;
        w1_rom[1558] = 2'b01;
        w1_rom[1559] = 2'b01;
        w1_rom[1560] = 2'b01;
        w1_rom[1561] = 2'b00;
        w1_rom[1562] = 2'b11;
        w1_rom[1563] = 2'b11;
        w1_rom[1564] = 2'b11;
        w1_rom[1565] = 2'b00;
        w1_rom[1566] = 2'b00;
        w1_rom[1567] = 2'b01;
        // Weights 1568-1583
        w1_rom[1568] = 2'b00;
        w1_rom[1569] = 2'b11;
        w1_rom[1570] = 2'b11;
        w1_rom[1571] = 2'b11;
        w1_rom[1572] = 2'b11;
        w1_rom[1573] = 2'b11;
        w1_rom[1574] = 2'b11;
        w1_rom[1575] = 2'b01;
        w1_rom[1576] = 2'b00;
        w1_rom[1577] = 2'b01;
        w1_rom[1578] = 2'b01;
        w1_rom[1579] = 2'b11;
        w1_rom[1580] = 2'b11;
        w1_rom[1581] = 2'b01;
        w1_rom[1582] = 2'b01;
        w1_rom[1583] = 2'b01;
        // Weights 1584-1599
        w1_rom[1584] = 2'b11;
        w1_rom[1585] = 2'b01;
        w1_rom[1586] = 2'b01;
        w1_rom[1587] = 2'b01;
        w1_rom[1588] = 2'b01;
        w1_rom[1589] = 2'b01;
        w1_rom[1590] = 2'b01;
        w1_rom[1591] = 2'b01;
        w1_rom[1592] = 2'b00;
        w1_rom[1593] = 2'b11;
        w1_rom[1594] = 2'b01;
        w1_rom[1595] = 2'b01;
        w1_rom[1596] = 2'b01;
        w1_rom[1597] = 2'b00;
        w1_rom[1598] = 2'b11;
        w1_rom[1599] = 2'b00;
        // Weights 1600-1615
        w1_rom[1600] = 2'b00;
        w1_rom[1601] = 2'b00;
        w1_rom[1602] = 2'b00;
        w1_rom[1603] = 2'b01;
        w1_rom[1604] = 2'b01;
        w1_rom[1605] = 2'b01;
        w1_rom[1606] = 2'b11;
        w1_rom[1607] = 2'b00;
        w1_rom[1608] = 2'b00;
        w1_rom[1609] = 2'b11;
        w1_rom[1610] = 2'b00;
        w1_rom[1611] = 2'b00;
        w1_rom[1612] = 2'b01;
        w1_rom[1613] = 2'b00;
        w1_rom[1614] = 2'b11;
        w1_rom[1615] = 2'b11;
        // Weights 1616-1631
        w1_rom[1616] = 2'b00;
        w1_rom[1617] = 2'b00;
        w1_rom[1618] = 2'b00;
        w1_rom[1619] = 2'b00;
        w1_rom[1620] = 2'b01;
        w1_rom[1621] = 2'b11;
        w1_rom[1622] = 2'b11;
        w1_rom[1623] = 2'b11;
        w1_rom[1624] = 2'b11;
        w1_rom[1625] = 2'b01;
        w1_rom[1626] = 2'b01;
        w1_rom[1627] = 2'b01;
        w1_rom[1628] = 2'b11;
        w1_rom[1629] = 2'b11;
        w1_rom[1630] = 2'b01;
        w1_rom[1631] = 2'b00;
        // Weights 1632-1647
        w1_rom[1632] = 2'b00;
        w1_rom[1633] = 2'b11;
        w1_rom[1634] = 2'b00;
        w1_rom[1635] = 2'b00;
        w1_rom[1636] = 2'b11;
        w1_rom[1637] = 2'b00;
        w1_rom[1638] = 2'b00;
        w1_rom[1639] = 2'b00;
        w1_rom[1640] = 2'b00;
        w1_rom[1641] = 2'b11;
        w1_rom[1642] = 2'b00;
        w1_rom[1643] = 2'b01;
        w1_rom[1644] = 2'b00;
        w1_rom[1645] = 2'b00;
        w1_rom[1646] = 2'b00;
        w1_rom[1647] = 2'b11;
        // Weights 1648-1663
        w1_rom[1648] = 2'b00;
        w1_rom[1649] = 2'b00;
        w1_rom[1650] = 2'b00;
        w1_rom[1651] = 2'b00;
        w1_rom[1652] = 2'b00;
        w1_rom[1653] = 2'b11;
        w1_rom[1654] = 2'b11;
        w1_rom[1655] = 2'b00;
        w1_rom[1656] = 2'b00;
        w1_rom[1657] = 2'b01;
        w1_rom[1658] = 2'b00;
        w1_rom[1659] = 2'b01;
        w1_rom[1660] = 2'b00;
        w1_rom[1661] = 2'b01;
        w1_rom[1662] = 2'b00;
        w1_rom[1663] = 2'b01;
        // Weights 1664-1679
        w1_rom[1664] = 2'b00;
        w1_rom[1665] = 2'b00;
        w1_rom[1666] = 2'b00;
        w1_rom[1667] = 2'b00;
        w1_rom[1668] = 2'b01;
        w1_rom[1669] = 2'b00;
        w1_rom[1670] = 2'b00;
        w1_rom[1671] = 2'b00;
        w1_rom[1672] = 2'b00;
        w1_rom[1673] = 2'b11;
        w1_rom[1674] = 2'b11;
        w1_rom[1675] = 2'b11;
        w1_rom[1676] = 2'b00;
        w1_rom[1677] = 2'b01;
        w1_rom[1678] = 2'b01;
        w1_rom[1679] = 2'b01;
        // Weights 1680-1695
        w1_rom[1680] = 2'b00;
        w1_rom[1681] = 2'b11;
        w1_rom[1682] = 2'b11;
        w1_rom[1683] = 2'b01;
        w1_rom[1684] = 2'b11;
        w1_rom[1685] = 2'b11;
        w1_rom[1686] = 2'b01;
        w1_rom[1687] = 2'b01;
        w1_rom[1688] = 2'b11;
        w1_rom[1689] = 2'b00;
        w1_rom[1690] = 2'b01;
        w1_rom[1691] = 2'b01;
        w1_rom[1692] = 2'b01;
        w1_rom[1693] = 2'b11;
        w1_rom[1694] = 2'b11;
        w1_rom[1695] = 2'b01;
        // Weights 1696-1711
        w1_rom[1696] = 2'b00;
        w1_rom[1697] = 2'b11;
        w1_rom[1698] = 2'b11;
        w1_rom[1699] = 2'b01;
        w1_rom[1700] = 2'b01;
        w1_rom[1701] = 2'b11;
        w1_rom[1702] = 2'b11;
        w1_rom[1703] = 2'b11;
        w1_rom[1704] = 2'b00;
        w1_rom[1705] = 2'b11;
        w1_rom[1706] = 2'b01;
        w1_rom[1707] = 2'b01;
        w1_rom[1708] = 2'b11;
        w1_rom[1709] = 2'b11;
        w1_rom[1710] = 2'b00;
        w1_rom[1711] = 2'b11;
        // Weights 1712-1727
        w1_rom[1712] = 2'b11;
        w1_rom[1713] = 2'b11;
        w1_rom[1714] = 2'b11;
        w1_rom[1715] = 2'b11;
        w1_rom[1716] = 2'b01;
        w1_rom[1717] = 2'b01;
        w1_rom[1718] = 2'b01;
        w1_rom[1719] = 2'b11;
        w1_rom[1720] = 2'b11;
        w1_rom[1721] = 2'b11;
        w1_rom[1722] = 2'b11;
        w1_rom[1723] = 2'b11;
        w1_rom[1724] = 2'b11;
        w1_rom[1725] = 2'b00;
        w1_rom[1726] = 2'b00;
        w1_rom[1727] = 2'b00;
        // Weights 1728-1743
        w1_rom[1728] = 2'b00;
        w1_rom[1729] = 2'b00;
        w1_rom[1730] = 2'b00;
        w1_rom[1731] = 2'b00;
        w1_rom[1732] = 2'b00;
        w1_rom[1733] = 2'b01;
        w1_rom[1734] = 2'b01;
        w1_rom[1735] = 2'b11;
        w1_rom[1736] = 2'b00;
        w1_rom[1737] = 2'b00;
        w1_rom[1738] = 2'b11;
        w1_rom[1739] = 2'b11;
        w1_rom[1740] = 2'b11;
        w1_rom[1741] = 2'b00;
        w1_rom[1742] = 2'b01;
        w1_rom[1743] = 2'b01;
        // Weights 1744-1759
        w1_rom[1744] = 2'b00;
        w1_rom[1745] = 2'b00;
        w1_rom[1746] = 2'b00;
        w1_rom[1747] = 2'b11;
        w1_rom[1748] = 2'b11;
        w1_rom[1749] = 2'b11;
        w1_rom[1750] = 2'b00;
        w1_rom[1751] = 2'b01;
        w1_rom[1752] = 2'b00;
        w1_rom[1753] = 2'b01;
        w1_rom[1754] = 2'b01;
        w1_rom[1755] = 2'b01;
        w1_rom[1756] = 2'b00;
        w1_rom[1757] = 2'b11;
        w1_rom[1758] = 2'b11;
        w1_rom[1759] = 2'b00;
        // Weights 1760-1775
        w1_rom[1760] = 2'b00;
        w1_rom[1761] = 2'b00;
        w1_rom[1762] = 2'b11;
        w1_rom[1763] = 2'b00;
        w1_rom[1764] = 2'b01;
        w1_rom[1765] = 2'b00;
        w1_rom[1766] = 2'b00;
        w1_rom[1767] = 2'b11;
        w1_rom[1768] = 2'b00;
        w1_rom[1769] = 2'b11;
        w1_rom[1770] = 2'b00;
        w1_rom[1771] = 2'b01;
        w1_rom[1772] = 2'b00;
        w1_rom[1773] = 2'b00;
        w1_rom[1774] = 2'b00;
        w1_rom[1775] = 2'b11;
        // Weights 1776-1791
        w1_rom[1776] = 2'b00;
        w1_rom[1777] = 2'b00;
        w1_rom[1778] = 2'b01;
        w1_rom[1779] = 2'b00;
        w1_rom[1780] = 2'b01;
        w1_rom[1781] = 2'b00;
        w1_rom[1782] = 2'b11;
        w1_rom[1783] = 2'b11;
        w1_rom[1784] = 2'b00;
        w1_rom[1785] = 2'b11;
        w1_rom[1786] = 2'b00;
        w1_rom[1787] = 2'b00;
        w1_rom[1788] = 2'b11;
        w1_rom[1789] = 2'b11;
        w1_rom[1790] = 2'b00;
        w1_rom[1791] = 2'b11;

        // Weights 1792-1807
        w1_rom[1792] = 2'b00;
        w1_rom[1793] = 2'b00;
        w1_rom[1794] = 2'b00;
        w1_rom[1795] = 2'b01;
        w1_rom[1796] = 2'b00;
        w1_rom[1797] = 2'b00;
        w1_rom[1798] = 2'b00;
        w1_rom[1799] = 2'b00;
        w1_rom[1800] = 2'b00;
        w1_rom[1801] = 2'b00;
        w1_rom[1802] = 2'b00;
        w1_rom[1803] = 2'b00;
        w1_rom[1804] = 2'b11;
        w1_rom[1805] = 2'b11;
        w1_rom[1806] = 2'b00;
        w1_rom[1807] = 2'b00;
        // Weights 1808-1823
        w1_rom[1808] = 2'b11;
        w1_rom[1809] = 2'b00;
        w1_rom[1810] = 2'b00;
        w1_rom[1811] = 2'b01;
        w1_rom[1812] = 2'b01;
        w1_rom[1813] = 2'b00;
        w1_rom[1814] = 2'b00;
        w1_rom[1815] = 2'b01;
        w1_rom[1816] = 2'b00;
        w1_rom[1817] = 2'b11;
        w1_rom[1818] = 2'b11;
        w1_rom[1819] = 2'b11;
        w1_rom[1820] = 2'b11;
        w1_rom[1821] = 2'b11;
        w1_rom[1822] = 2'b11;
        w1_rom[1823] = 2'b00;
        // Weights 1824-1839
        w1_rom[1824] = 2'b00;
        w1_rom[1825] = 2'b00;
        w1_rom[1826] = 2'b00;
        w1_rom[1827] = 2'b11;
        w1_rom[1828] = 2'b00;
        w1_rom[1829] = 2'b00;
        w1_rom[1830] = 2'b11;
        w1_rom[1831] = 2'b01;
        w1_rom[1832] = 2'b00;
        w1_rom[1833] = 2'b01;
        w1_rom[1834] = 2'b11;
        w1_rom[1835] = 2'b01;
        w1_rom[1836] = 2'b00;
        w1_rom[1837] = 2'b00;
        w1_rom[1838] = 2'b00;
        w1_rom[1839] = 2'b01;
        // Weights 1840-1855
        w1_rom[1840] = 2'b00;
        w1_rom[1841] = 2'b00;
        w1_rom[1842] = 2'b00;
        w1_rom[1843] = 2'b00;
        w1_rom[1844] = 2'b11;
        w1_rom[1845] = 2'b00;
        w1_rom[1846] = 2'b01;
        w1_rom[1847] = 2'b01;
        w1_rom[1848] = 2'b00;
        w1_rom[1849] = 2'b00;
        w1_rom[1850] = 2'b11;
        w1_rom[1851] = 2'b00;
        w1_rom[1852] = 2'b01;
        w1_rom[1853] = 2'b00;
        w1_rom[1854] = 2'b11;
        w1_rom[1855] = 2'b00;
        // Weights 1856-1871
        w1_rom[1856] = 2'b01;
        w1_rom[1857] = 2'b01;
        w1_rom[1858] = 2'b00;
        w1_rom[1859] = 2'b00;
        w1_rom[1860] = 2'b00;
        w1_rom[1861] = 2'b00;
        w1_rom[1862] = 2'b00;
        w1_rom[1863] = 2'b00;
        w1_rom[1864] = 2'b00;
        w1_rom[1865] = 2'b00;
        w1_rom[1866] = 2'b01;
        w1_rom[1867] = 2'b00;
        w1_rom[1868] = 2'b00;
        w1_rom[1869] = 2'b00;
        w1_rom[1870] = 2'b00;
        w1_rom[1871] = 2'b01;
        // Weights 1872-1887
        w1_rom[1872] = 2'b00;
        w1_rom[1873] = 2'b01;
        w1_rom[1874] = 2'b01;
        w1_rom[1875] = 2'b11;
        w1_rom[1876] = 2'b11;
        w1_rom[1877] = 2'b00;
        w1_rom[1878] = 2'b00;
        w1_rom[1879] = 2'b11;
        w1_rom[1880] = 2'b00;
        w1_rom[1881] = 2'b11;
        w1_rom[1882] = 2'b11;
        w1_rom[1883] = 2'b11;
        w1_rom[1884] = 2'b11;
        w1_rom[1885] = 2'b01;
        w1_rom[1886] = 2'b11;
        w1_rom[1887] = 2'b11;
        // Weights 1888-1903
        w1_rom[1888] = 2'b00;
        w1_rom[1889] = 2'b00;
        w1_rom[1890] = 2'b01;
        w1_rom[1891] = 2'b01;
        w1_rom[1892] = 2'b01;
        w1_rom[1893] = 2'b01;
        w1_rom[1894] = 2'b00;
        w1_rom[1895] = 2'b01;
        w1_rom[1896] = 2'b01;
        w1_rom[1897] = 2'b01;
        w1_rom[1898] = 2'b01;
        w1_rom[1899] = 2'b01;
        w1_rom[1900] = 2'b01;
        w1_rom[1901] = 2'b01;
        w1_rom[1902] = 2'b01;
        w1_rom[1903] = 2'b01;
        // Weights 1904-1919
        w1_rom[1904] = 2'b00;
        w1_rom[1905] = 2'b00;
        w1_rom[1906] = 2'b11;
        w1_rom[1907] = 2'b11;
        w1_rom[1908] = 2'b11;
        w1_rom[1909] = 2'b01;
        w1_rom[1910] = 2'b01;
        w1_rom[1911] = 2'b01;
        w1_rom[1912] = 2'b00;
        w1_rom[1913] = 2'b11;
        w1_rom[1914] = 2'b00;
        w1_rom[1915] = 2'b11;
        w1_rom[1916] = 2'b11;
        w1_rom[1917] = 2'b11;
        w1_rom[1918] = 2'b11;
        w1_rom[1919] = 2'b00;
        // Weights 1920-1935
        w1_rom[1920] = 2'b11;
        w1_rom[1921] = 2'b00;
        w1_rom[1922] = 2'b00;
        w1_rom[1923] = 2'b11;
        w1_rom[1924] = 2'b01;
        w1_rom[1925] = 2'b00;
        w1_rom[1926] = 2'b00;
        w1_rom[1927] = 2'b01;
        w1_rom[1928] = 2'b01;
        w1_rom[1929] = 2'b01;
        w1_rom[1930] = 2'b01;
        w1_rom[1931] = 2'b00;
        w1_rom[1932] = 2'b00;
        w1_rom[1933] = 2'b01;
        w1_rom[1934] = 2'b11;
        w1_rom[1935] = 2'b00;
        // Weights 1936-1951
        w1_rom[1936] = 2'b00;
        w1_rom[1937] = 2'b00;
        w1_rom[1938] = 2'b11;
        w1_rom[1939] = 2'b00;
        w1_rom[1940] = 2'b01;
        w1_rom[1941] = 2'b00;
        w1_rom[1942] = 2'b00;
        w1_rom[1943] = 2'b11;
        w1_rom[1944] = 2'b00;
        w1_rom[1945] = 2'b11;
        w1_rom[1946] = 2'b00;
        w1_rom[1947] = 2'b11;
        w1_rom[1948] = 2'b01;
        w1_rom[1949] = 2'b01;
        w1_rom[1950] = 2'b00;
        w1_rom[1951] = 2'b11;
        // Weights 1952-1967
        w1_rom[1952] = 2'b01;
        w1_rom[1953] = 2'b01;
        w1_rom[1954] = 2'b01;
        w1_rom[1955] = 2'b00;
        w1_rom[1956] = 2'b00;
        w1_rom[1957] = 2'b00;
        w1_rom[1958] = 2'b01;
        w1_rom[1959] = 2'b11;
        w1_rom[1960] = 2'b00;
        w1_rom[1961] = 2'b11;
        w1_rom[1962] = 2'b00;
        w1_rom[1963] = 2'b11;
        w1_rom[1964] = 2'b00;
        w1_rom[1965] = 2'b01;
        w1_rom[1966] = 2'b11;
        w1_rom[1967] = 2'b11;
        // Weights 1968-1983
        w1_rom[1968] = 2'b01;
        w1_rom[1969] = 2'b01;
        w1_rom[1970] = 2'b11;
        w1_rom[1971] = 2'b11;
        w1_rom[1972] = 2'b00;
        w1_rom[1973] = 2'b00;
        w1_rom[1974] = 2'b11;
        w1_rom[1975] = 2'b11;
        w1_rom[1976] = 2'b00;
        w1_rom[1977] = 2'b01;
        w1_rom[1978] = 2'b01;
        w1_rom[1979] = 2'b11;
        w1_rom[1980] = 2'b11;
        w1_rom[1981] = 2'b11;
        w1_rom[1982] = 2'b01;
        w1_rom[1983] = 2'b00;
        // Weights 1984-1999
        w1_rom[1984] = 2'b00;
        w1_rom[1985] = 2'b00;
        w1_rom[1986] = 2'b00;
        w1_rom[1987] = 2'b11;
        w1_rom[1988] = 2'b00;
        w1_rom[1989] = 2'b11;
        w1_rom[1990] = 2'b00;
        w1_rom[1991] = 2'b00;
        w1_rom[1992] = 2'b00;
        w1_rom[1993] = 2'b00;
        w1_rom[1994] = 2'b00;
        w1_rom[1995] = 2'b11;
        w1_rom[1996] = 2'b11;
        w1_rom[1997] = 2'b00;
        w1_rom[1998] = 2'b00;
        w1_rom[1999] = 2'b00;
        // Weights 2000-2015
        w1_rom[2000] = 2'b01;
        w1_rom[2001] = 2'b01;
        w1_rom[2002] = 2'b00;
        w1_rom[2003] = 2'b00;
        w1_rom[2004] = 2'b11;
        w1_rom[2005] = 2'b00;
        w1_rom[2006] = 2'b01;
        w1_rom[2007] = 2'b01;
        w1_rom[2008] = 2'b00;
        w1_rom[2009] = 2'b01;
        w1_rom[2010] = 2'b00;
        w1_rom[2011] = 2'b01;
        w1_rom[2012] = 2'b01;
        w1_rom[2013] = 2'b11;
        w1_rom[2014] = 2'b11;
        w1_rom[2015] = 2'b00;
        // Weights 2016-2031
        w1_rom[2016] = 2'b00;
        w1_rom[2017] = 2'b00;
        w1_rom[2018] = 2'b00;
        w1_rom[2019] = 2'b00;
        w1_rom[2020] = 2'b00;
        w1_rom[2021] = 2'b01;
        w1_rom[2022] = 2'b00;
        w1_rom[2023] = 2'b00;
        w1_rom[2024] = 2'b00;
        w1_rom[2025] = 2'b00;
        w1_rom[2026] = 2'b00;
        w1_rom[2027] = 2'b11;
        w1_rom[2028] = 2'b00;
        w1_rom[2029] = 2'b00;
        w1_rom[2030] = 2'b00;
        w1_rom[2031] = 2'b11;
        // Weights 2032-2047
        w1_rom[2032] = 2'b01;
        w1_rom[2033] = 2'b00;
        w1_rom[2034] = 2'b00;
        w1_rom[2035] = 2'b00;
        w1_rom[2036] = 2'b00;
        w1_rom[2037] = 2'b00;
        w1_rom[2038] = 2'b11;
        w1_rom[2039] = 2'b00;
        w1_rom[2040] = 2'b00;
        w1_rom[2041] = 2'b01;
        w1_rom[2042] = 2'b01;
        w1_rom[2043] = 2'b00;
        w1_rom[2044] = 2'b00;
        w1_rom[2045] = 2'b11;
        w1_rom[2046] = 2'b00;
        w1_rom[2047] = 2'b00;

        // Weights 2048-2063
        w1_rom[2048] = 2'b00;
        w1_rom[2049] = 2'b00;
        w1_rom[2050] = 2'b00;
        w1_rom[2051] = 2'b11;
        w1_rom[2052] = 2'b00;
        w1_rom[2053] = 2'b00;
        w1_rom[2054] = 2'b00;
        w1_rom[2055] = 2'b00;
        w1_rom[2056] = 2'b00;
        w1_rom[2057] = 2'b00;
        w1_rom[2058] = 2'b00;
        w1_rom[2059] = 2'b00;
        w1_rom[2060] = 2'b00;
        w1_rom[2061] = 2'b00;
        w1_rom[2062] = 2'b00;
        w1_rom[2063] = 2'b11;
        // Weights 2064-2079
        w1_rom[2064] = 2'b00;
        w1_rom[2065] = 2'b01;
        w1_rom[2066] = 2'b01;
        w1_rom[2067] = 2'b00;
        w1_rom[2068] = 2'b11;
        w1_rom[2069] = 2'b01;
        w1_rom[2070] = 2'b01;
        w1_rom[2071] = 2'b11;
        w1_rom[2072] = 2'b01;
        w1_rom[2073] = 2'b11;
        w1_rom[2074] = 2'b11;
        w1_rom[2075] = 2'b11;
        w1_rom[2076] = 2'b00;
        w1_rom[2077] = 2'b01;
        w1_rom[2078] = 2'b01;
        w1_rom[2079] = 2'b00;
        // Weights 2080-2095
        w1_rom[2080] = 2'b11;
        w1_rom[2081] = 2'b11;
        w1_rom[2082] = 2'b11;
        w1_rom[2083] = 2'b01;
        w1_rom[2084] = 2'b01;
        w1_rom[2085] = 2'b11;
        w1_rom[2086] = 2'b11;
        w1_rom[2087] = 2'b01;
        w1_rom[2088] = 2'b00;
        w1_rom[2089] = 2'b00;
        w1_rom[2090] = 2'b01;
        w1_rom[2091] = 2'b01;
        w1_rom[2092] = 2'b00;
        w1_rom[2093] = 2'b11;
        w1_rom[2094] = 2'b00;
        w1_rom[2095] = 2'b01;
        // Weights 2096-2111
        w1_rom[2096] = 2'b01;
        w1_rom[2097] = 2'b01;
        w1_rom[2098] = 2'b00;
        w1_rom[2099] = 2'b11;
        w1_rom[2100] = 2'b01;
        w1_rom[2101] = 2'b01;
        w1_rom[2102] = 2'b01;
        w1_rom[2103] = 2'b01;
        w1_rom[2104] = 2'b11;
        w1_rom[2105] = 2'b11;
        w1_rom[2106] = 2'b11;
        w1_rom[2107] = 2'b11;
        w1_rom[2108] = 2'b00;
        w1_rom[2109] = 2'b11;
        w1_rom[2110] = 2'b11;
        w1_rom[2111] = 2'b01;
        // Weights 2112-2127
        w1_rom[2112] = 2'b11;
        w1_rom[2113] = 2'b00;
        w1_rom[2114] = 2'b11;
        w1_rom[2115] = 2'b00;
        w1_rom[2116] = 2'b00;
        w1_rom[2117] = 2'b00;
        w1_rom[2118] = 2'b11;
        w1_rom[2119] = 2'b00;
        w1_rom[2120] = 2'b00;
        w1_rom[2121] = 2'b00;
        w1_rom[2122] = 2'b00;
        w1_rom[2123] = 2'b00;
        w1_rom[2124] = 2'b00;
        w1_rom[2125] = 2'b00;
        w1_rom[2126] = 2'b00;
        w1_rom[2127] = 2'b11;
        // Weights 2128-2143
        w1_rom[2128] = 2'b00;
        w1_rom[2129] = 2'b01;
        w1_rom[2130] = 2'b00;
        w1_rom[2131] = 2'b11;
        w1_rom[2132] = 2'b00;
        w1_rom[2133] = 2'b00;
        w1_rom[2134] = 2'b11;
        w1_rom[2135] = 2'b11;
        w1_rom[2136] = 2'b11;
        w1_rom[2137] = 2'b00;
        w1_rom[2138] = 2'b11;
        w1_rom[2139] = 2'b11;
        w1_rom[2140] = 2'b00;
        w1_rom[2141] = 2'b01;
        w1_rom[2142] = 2'b01;
        w1_rom[2143] = 2'b11;
        // Weights 2144-2159
        w1_rom[2144] = 2'b00;
        w1_rom[2145] = 2'b01;
        w1_rom[2146] = 2'b00;
        w1_rom[2147] = 2'b00;
        w1_rom[2148] = 2'b00;
        w1_rom[2149] = 2'b00;
        w1_rom[2150] = 2'b01;
        w1_rom[2151] = 2'b00;
        w1_rom[2152] = 2'b00;
        w1_rom[2153] = 2'b11;
        w1_rom[2154] = 2'b01;
        w1_rom[2155] = 2'b01;
        w1_rom[2156] = 2'b00;
        w1_rom[2157] = 2'b11;
        w1_rom[2158] = 2'b11;
        w1_rom[2159] = 2'b00;
        // Weights 2160-2175
        w1_rom[2160] = 2'b00;
        w1_rom[2161] = 2'b00;
        w1_rom[2162] = 2'b11;
        w1_rom[2163] = 2'b01;
        w1_rom[2164] = 2'b01;
        w1_rom[2165] = 2'b00;
        w1_rom[2166] = 2'b00;
        w1_rom[2167] = 2'b00;
        w1_rom[2168] = 2'b00;
        w1_rom[2169] = 2'b00;
        w1_rom[2170] = 2'b11;
        w1_rom[2171] = 2'b11;
        w1_rom[2172] = 2'b11;
        w1_rom[2173] = 2'b00;
        w1_rom[2174] = 2'b11;
        w1_rom[2175] = 2'b00;
        // Weights 2176-2191
        w1_rom[2176] = 2'b01;
        w1_rom[2177] = 2'b00;
        w1_rom[2178] = 2'b00;
        w1_rom[2179] = 2'b01;
        w1_rom[2180] = 2'b01;
        w1_rom[2181] = 2'b01;
        w1_rom[2182] = 2'b01;
        w1_rom[2183] = 2'b11;
        w1_rom[2184] = 2'b01;
        w1_rom[2185] = 2'b11;
        w1_rom[2186] = 2'b01;
        w1_rom[2187] = 2'b11;
        w1_rom[2188] = 2'b11;
        w1_rom[2189] = 2'b00;
        w1_rom[2190] = 2'b01;
        w1_rom[2191] = 2'b01;
        // Weights 2192-2207
        w1_rom[2192] = 2'b00;
        w1_rom[2193] = 2'b01;
        w1_rom[2194] = 2'b01;
        w1_rom[2195] = 2'b11;
        w1_rom[2196] = 2'b11;
        w1_rom[2197] = 2'b11;
        w1_rom[2198] = 2'b01;
        w1_rom[2199] = 2'b01;
        w1_rom[2200] = 2'b01;
        w1_rom[2201] = 2'b00;
        w1_rom[2202] = 2'b01;
        w1_rom[2203] = 2'b01;
        w1_rom[2204] = 2'b11;
        w1_rom[2205] = 2'b11;
        w1_rom[2206] = 2'b11;
        w1_rom[2207] = 2'b01;
        // Weights 2208-2223
        w1_rom[2208] = 2'b00;
        w1_rom[2209] = 2'b11;
        w1_rom[2210] = 2'b11;
        w1_rom[2211] = 2'b11;
        w1_rom[2212] = 2'b11;
        w1_rom[2213] = 2'b01;
        w1_rom[2214] = 2'b01;
        w1_rom[2215] = 2'b01;
        w1_rom[2216] = 2'b00;
        w1_rom[2217] = 2'b01;
        w1_rom[2218] = 2'b01;
        w1_rom[2219] = 2'b01;
        w1_rom[2220] = 2'b00;
        w1_rom[2221] = 2'b01;
        w1_rom[2222] = 2'b01;
        w1_rom[2223] = 2'b00;
        // Weights 2224-2239
        w1_rom[2224] = 2'b00;
        w1_rom[2225] = 2'b11;
        w1_rom[2226] = 2'b00;
        w1_rom[2227] = 2'b01;
        w1_rom[2228] = 2'b00;
        w1_rom[2229] = 2'b11;
        w1_rom[2230] = 2'b11;
        w1_rom[2231] = 2'b00;
        w1_rom[2232] = 2'b11;
        w1_rom[2233] = 2'b00;
        w1_rom[2234] = 2'b11;
        w1_rom[2235] = 2'b01;
        w1_rom[2236] = 2'b00;
        w1_rom[2237] = 2'b11;
        w1_rom[2238] = 2'b11;
        w1_rom[2239] = 2'b00;
        // Weights 2240-2255
        w1_rom[2240] = 2'b00;
        w1_rom[2241] = 2'b00;
        w1_rom[2242] = 2'b11;
        w1_rom[2243] = 2'b11;
        w1_rom[2244] = 2'b11;
        w1_rom[2245] = 2'b11;
        w1_rom[2246] = 2'b11;
        w1_rom[2247] = 2'b00;
        w1_rom[2248] = 2'b00;
        w1_rom[2249] = 2'b00;
        w1_rom[2250] = 2'b11;
        w1_rom[2251] = 2'b11;
        w1_rom[2252] = 2'b11;
        w1_rom[2253] = 2'b11;
        w1_rom[2254] = 2'b01;
        w1_rom[2255] = 2'b00;
        // Weights 2256-2271
        w1_rom[2256] = 2'b00;
        w1_rom[2257] = 2'b11;
        w1_rom[2258] = 2'b00;
        w1_rom[2259] = 2'b01;
        w1_rom[2260] = 2'b00;
        w1_rom[2261] = 2'b01;
        w1_rom[2262] = 2'b01;
        w1_rom[2263] = 2'b11;
        w1_rom[2264] = 2'b01;
        w1_rom[2265] = 2'b01;
        w1_rom[2266] = 2'b01;
        w1_rom[2267] = 2'b11;
        w1_rom[2268] = 2'b11;
        w1_rom[2269] = 2'b01;
        w1_rom[2270] = 2'b11;
        w1_rom[2271] = 2'b11;
        // Weights 2272-2287
        w1_rom[2272] = 2'b00;
        w1_rom[2273] = 2'b01;
        w1_rom[2274] = 2'b01;
        w1_rom[2275] = 2'b11;
        w1_rom[2276] = 2'b01;
        w1_rom[2277] = 2'b01;
        w1_rom[2278] = 2'b11;
        w1_rom[2279] = 2'b11;
        w1_rom[2280] = 2'b11;
        w1_rom[2281] = 2'b11;
        w1_rom[2282] = 2'b11;
        w1_rom[2283] = 2'b11;
        w1_rom[2284] = 2'b01;
        w1_rom[2285] = 2'b11;
        w1_rom[2286] = 2'b11;
        w1_rom[2287] = 2'b01;
        // Weights 2288-2303
        w1_rom[2288] = 2'b11;
        w1_rom[2289] = 2'b11;
        w1_rom[2290] = 2'b11;
        w1_rom[2291] = 2'b11;
        w1_rom[2292] = 2'b11;
        w1_rom[2293] = 2'b01;
        w1_rom[2294] = 2'b01;
        w1_rom[2295] = 2'b01;
        w1_rom[2296] = 2'b01;
        w1_rom[2297] = 2'b01;
        w1_rom[2298] = 2'b01;
        w1_rom[2299] = 2'b01;
        w1_rom[2300] = 2'b01;
        w1_rom[2301] = 2'b01;
        w1_rom[2302] = 2'b01;
        w1_rom[2303] = 2'b00;

        // Weights 2304-2319
        w1_rom[2304] = 2'b00;
        w1_rom[2305] = 2'b00;
        w1_rom[2306] = 2'b00;
        w1_rom[2307] = 2'b00;
        w1_rom[2308] = 2'b00;
        w1_rom[2309] = 2'b00;
        w1_rom[2310] = 2'b00;
        w1_rom[2311] = 2'b11;
        w1_rom[2312] = 2'b00;
        w1_rom[2313] = 2'b00;
        w1_rom[2314] = 2'b00;
        w1_rom[2315] = 2'b11;
        w1_rom[2316] = 2'b11;
        w1_rom[2317] = 2'b11;
        w1_rom[2318] = 2'b01;
        w1_rom[2319] = 2'b01;
        // Weights 2320-2335
        w1_rom[2320] = 2'b00;
        w1_rom[2321] = 2'b01;
        w1_rom[2322] = 2'b01;
        w1_rom[2323] = 2'b00;
        w1_rom[2324] = 2'b11;
        w1_rom[2325] = 2'b00;
        w1_rom[2326] = 2'b01;
        w1_rom[2327] = 2'b01;
        w1_rom[2328] = 2'b01;
        w1_rom[2329] = 2'b01;
        w1_rom[2330] = 2'b01;
        w1_rom[2331] = 2'b01;
        w1_rom[2332] = 2'b01;
        w1_rom[2333] = 2'b01;
        w1_rom[2334] = 2'b11;
        w1_rom[2335] = 2'b11;
        // Weights 2336-2351
        w1_rom[2336] = 2'b00;
        w1_rom[2337] = 2'b11;
        w1_rom[2338] = 2'b11;
        w1_rom[2339] = 2'b11;
        w1_rom[2340] = 2'b01;
        w1_rom[2341] = 2'b01;
        w1_rom[2342] = 2'b01;
        w1_rom[2343] = 2'b11;
        w1_rom[2344] = 2'b00;
        w1_rom[2345] = 2'b00;
        w1_rom[2346] = 2'b11;
        w1_rom[2347] = 2'b11;
        w1_rom[2348] = 2'b00;
        w1_rom[2349] = 2'b11;
        w1_rom[2350] = 2'b11;
        w1_rom[2351] = 2'b11;
        // Weights 2352-2367
        w1_rom[2352] = 2'b00;
        w1_rom[2353] = 2'b00;
        w1_rom[2354] = 2'b00;
        w1_rom[2355] = 2'b01;
        w1_rom[2356] = 2'b00;
        w1_rom[2357] = 2'b11;
        w1_rom[2358] = 2'b11;
        w1_rom[2359] = 2'b00;
        w1_rom[2360] = 2'b11;
        w1_rom[2361] = 2'b01;
        w1_rom[2362] = 2'b01;
        w1_rom[2363] = 2'b01;
        w1_rom[2364] = 2'b01;
        w1_rom[2365] = 2'b00;
        w1_rom[2366] = 2'b11;
        w1_rom[2367] = 2'b00;
        // Weights 2368-2383
        w1_rom[2368] = 2'b00;
        w1_rom[2369] = 2'b00;
        w1_rom[2370] = 2'b00;
        w1_rom[2371] = 2'b00;
        w1_rom[2372] = 2'b00;
        w1_rom[2373] = 2'b00;
        w1_rom[2374] = 2'b00;
        w1_rom[2375] = 2'b01;
        w1_rom[2376] = 2'b00;
        w1_rom[2377] = 2'b01;
        w1_rom[2378] = 2'b01;
        w1_rom[2379] = 2'b00;
        w1_rom[2380] = 2'b01;
        w1_rom[2381] = 2'b00;
        w1_rom[2382] = 2'b11;
        w1_rom[2383] = 2'b00;
        // Weights 2384-2399
        w1_rom[2384] = 2'b00;
        w1_rom[2385] = 2'b01;
        w1_rom[2386] = 2'b00;
        w1_rom[2387] = 2'b01;
        w1_rom[2388] = 2'b01;
        w1_rom[2389] = 2'b01;
        w1_rom[2390] = 2'b00;
        w1_rom[2391] = 2'b00;
        w1_rom[2392] = 2'b00;
        w1_rom[2393] = 2'b11;
        w1_rom[2394] = 2'b11;
        w1_rom[2395] = 2'b11;
        w1_rom[2396] = 2'b00;
        w1_rom[2397] = 2'b01;
        w1_rom[2398] = 2'b00;
        w1_rom[2399] = 2'b00;
        // Weights 2400-2415
        w1_rom[2400] = 2'b11;
        w1_rom[2401] = 2'b01;
        w1_rom[2402] = 2'b00;
        w1_rom[2403] = 2'b11;
        w1_rom[2404] = 2'b00;
        w1_rom[2405] = 2'b11;
        w1_rom[2406] = 2'b00;
        w1_rom[2407] = 2'b00;
        w1_rom[2408] = 2'b00;
        w1_rom[2409] = 2'b01;
        w1_rom[2410] = 2'b00;
        w1_rom[2411] = 2'b11;
        w1_rom[2412] = 2'b00;
        w1_rom[2413] = 2'b00;
        w1_rom[2414] = 2'b00;
        w1_rom[2415] = 2'b00;
        // Weights 2416-2431
        w1_rom[2416] = 2'b00;
        w1_rom[2417] = 2'b00;
        w1_rom[2418] = 2'b11;
        w1_rom[2419] = 2'b11;
        w1_rom[2420] = 2'b11;
        w1_rom[2421] = 2'b11;
        w1_rom[2422] = 2'b00;
        w1_rom[2423] = 2'b00;
        w1_rom[2424] = 2'b00;
        w1_rom[2425] = 2'b00;
        w1_rom[2426] = 2'b01;
        w1_rom[2427] = 2'b01;
        w1_rom[2428] = 2'b00;
        w1_rom[2429] = 2'b00;
        w1_rom[2430] = 2'b00;
        w1_rom[2431] = 2'b00;
        // Weights 2432-2447
        w1_rom[2432] = 2'b00;
        w1_rom[2433] = 2'b01;
        w1_rom[2434] = 2'b01;
        w1_rom[2435] = 2'b01;
        w1_rom[2436] = 2'b01;
        w1_rom[2437] = 2'b01;
        w1_rom[2438] = 2'b00;
        w1_rom[2439] = 2'b11;
        w1_rom[2440] = 2'b00;
        w1_rom[2441] = 2'b00;
        w1_rom[2442] = 2'b00;
        w1_rom[2443] = 2'b11;
        w1_rom[2444] = 2'b11;
        w1_rom[2445] = 2'b00;
        w1_rom[2446] = 2'b01;
        w1_rom[2447] = 2'b01;
        // Weights 2448-2463
        w1_rom[2448] = 2'b00;
        w1_rom[2449] = 2'b00;
        w1_rom[2450] = 2'b01;
        w1_rom[2451] = 2'b11;
        w1_rom[2452] = 2'b11;
        w1_rom[2453] = 2'b11;
        w1_rom[2454] = 2'b00;
        w1_rom[2455] = 2'b01;
        w1_rom[2456] = 2'b00;
        w1_rom[2457] = 2'b00;
        w1_rom[2458] = 2'b00;
        w1_rom[2459] = 2'b01;
        w1_rom[2460] = 2'b01;
        w1_rom[2461] = 2'b11;
        w1_rom[2462] = 2'b11;
        w1_rom[2463] = 2'b00;
        // Weights 2464-2479
        w1_rom[2464] = 2'b00;
        w1_rom[2465] = 2'b11;
        w1_rom[2466] = 2'b00;
        w1_rom[2467] = 2'b11;
        w1_rom[2468] = 2'b01;
        w1_rom[2469] = 2'b01;
        w1_rom[2470] = 2'b01;
        w1_rom[2471] = 2'b00;
        w1_rom[2472] = 2'b00;
        w1_rom[2473] = 2'b11;
        w1_rom[2474] = 2'b11;
        w1_rom[2475] = 2'b00;
        w1_rom[2476] = 2'b00;
        w1_rom[2477] = 2'b01;
        w1_rom[2478] = 2'b00;
        w1_rom[2479] = 2'b11;
        // Weights 2480-2495
        w1_rom[2480] = 2'b00;
        w1_rom[2481] = 2'b11;
        w1_rom[2482] = 2'b00;
        w1_rom[2483] = 2'b01;
        w1_rom[2484] = 2'b00;
        w1_rom[2485] = 2'b00;
        w1_rom[2486] = 2'b11;
        w1_rom[2487] = 2'b11;
        w1_rom[2488] = 2'b01;
        w1_rom[2489] = 2'b00;
        w1_rom[2490] = 2'b01;
        w1_rom[2491] = 2'b00;
        w1_rom[2492] = 2'b00;
        w1_rom[2493] = 2'b11;
        w1_rom[2494] = 2'b00;
        w1_rom[2495] = 2'b00;
        // Weights 2496-2511
        w1_rom[2496] = 2'b11;
        w1_rom[2497] = 2'b00;
        w1_rom[2498] = 2'b01;
        w1_rom[2499] = 2'b11;
        w1_rom[2500] = 2'b00;
        w1_rom[2501] = 2'b11;
        w1_rom[2502] = 2'b00;
        w1_rom[2503] = 2'b00;
        w1_rom[2504] = 2'b00;
        w1_rom[2505] = 2'b00;
        w1_rom[2506] = 2'b00;
        w1_rom[2507] = 2'b01;
        w1_rom[2508] = 2'b00;
        w1_rom[2509] = 2'b00;
        w1_rom[2510] = 2'b00;
        w1_rom[2511] = 2'b01;
        // Weights 2512-2527
        w1_rom[2512] = 2'b01;
        w1_rom[2513] = 2'b01;
        w1_rom[2514] = 2'b00;
        w1_rom[2515] = 2'b01;
        w1_rom[2516] = 2'b00;
        w1_rom[2517] = 2'b01;
        w1_rom[2518] = 2'b01;
        w1_rom[2519] = 2'b01;
        w1_rom[2520] = 2'b01;
        w1_rom[2521] = 2'b00;
        w1_rom[2522] = 2'b00;
        w1_rom[2523] = 2'b11;
        w1_rom[2524] = 2'b01;
        w1_rom[2525] = 2'b00;
        w1_rom[2526] = 2'b11;
        w1_rom[2527] = 2'b01;
        // Weights 2528-2543
        w1_rom[2528] = 2'b11;
        w1_rom[2529] = 2'b11;
        w1_rom[2530] = 2'b11;
        w1_rom[2531] = 2'b11;
        w1_rom[2532] = 2'b01;
        w1_rom[2533] = 2'b00;
        w1_rom[2534] = 2'b11;
        w1_rom[2535] = 2'b00;
        w1_rom[2536] = 2'b00;
        w1_rom[2537] = 2'b01;
        w1_rom[2538] = 2'b00;
        w1_rom[2539] = 2'b11;
        w1_rom[2540] = 2'b00;
        w1_rom[2541] = 2'b11;
        w1_rom[2542] = 2'b00;
        w1_rom[2543] = 2'b01;
        // Weights 2544-2559
        w1_rom[2544] = 2'b00;
        w1_rom[2545] = 2'b00;
        w1_rom[2546] = 2'b01;
        w1_rom[2547] = 2'b11;
        w1_rom[2548] = 2'b00;
        w1_rom[2549] = 2'b01;
        w1_rom[2550] = 2'b01;
        w1_rom[2551] = 2'b00;
        w1_rom[2552] = 2'b00;
        w1_rom[2553] = 2'b11;
        w1_rom[2554] = 2'b11;
        w1_rom[2555] = 2'b01;
        w1_rom[2556] = 2'b00;
        w1_rom[2557] = 2'b01;
        w1_rom[2558] = 2'b00;
        w1_rom[2559] = 2'b00;

        // Weights 2560-2575
        w1_rom[2560] = 2'b00;
        w1_rom[2561] = 2'b00;
        w1_rom[2562] = 2'b00;
        w1_rom[2563] = 2'b11;
        w1_rom[2564] = 2'b00;
        w1_rom[2565] = 2'b00;
        w1_rom[2566] = 2'b11;
        w1_rom[2567] = 2'b01;
        w1_rom[2568] = 2'b11;
        w1_rom[2569] = 2'b11;
        w1_rom[2570] = 2'b00;
        w1_rom[2571] = 2'b11;
        w1_rom[2572] = 2'b11;
        w1_rom[2573] = 2'b00;
        w1_rom[2574] = 2'b01;
        w1_rom[2575] = 2'b01;
        // Weights 2576-2591
        w1_rom[2576] = 2'b00;
        w1_rom[2577] = 2'b00;
        w1_rom[2578] = 2'b01;
        w1_rom[2579] = 2'b00;
        w1_rom[2580] = 2'b11;
        w1_rom[2581] = 2'b00;
        w1_rom[2582] = 2'b01;
        w1_rom[2583] = 2'b01;
        w1_rom[2584] = 2'b00;
        w1_rom[2585] = 2'b01;
        w1_rom[2586] = 2'b01;
        w1_rom[2587] = 2'b01;
        w1_rom[2588] = 2'b11;
        w1_rom[2589] = 2'b11;
        w1_rom[2590] = 2'b00;
        w1_rom[2591] = 2'b00;
        // Weights 2592-2607
        w1_rom[2592] = 2'b00;
        w1_rom[2593] = 2'b00;
        w1_rom[2594] = 2'b11;
        w1_rom[2595] = 2'b00;
        w1_rom[2596] = 2'b00;
        w1_rom[2597] = 2'b00;
        w1_rom[2598] = 2'b01;
        w1_rom[2599] = 2'b11;
        w1_rom[2600] = 2'b00;
        w1_rom[2601] = 2'b11;
        w1_rom[2602] = 2'b00;
        w1_rom[2603] = 2'b01;
        w1_rom[2604] = 2'b00;
        w1_rom[2605] = 2'b00;
        w1_rom[2606] = 2'b00;
        w1_rom[2607] = 2'b00;
        // Weights 2608-2623
        w1_rom[2608] = 2'b11;
        w1_rom[2609] = 2'b11;
        w1_rom[2610] = 2'b00;
        w1_rom[2611] = 2'b01;
        w1_rom[2612] = 2'b01;
        w1_rom[2613] = 2'b11;
        w1_rom[2614] = 2'b00;
        w1_rom[2615] = 2'b00;
        w1_rom[2616] = 2'b00;
        w1_rom[2617] = 2'b11;
        w1_rom[2618] = 2'b11;
        w1_rom[2619] = 2'b00;
        w1_rom[2620] = 2'b00;
        w1_rom[2621] = 2'b00;
        w1_rom[2622] = 2'b00;
        w1_rom[2623] = 2'b00;
        // Weights 2624-2639
        w1_rom[2624] = 2'b00;
        w1_rom[2625] = 2'b00;
        w1_rom[2626] = 2'b00;
        w1_rom[2627] = 2'b00;
        w1_rom[2628] = 2'b01;
        w1_rom[2629] = 2'b01;
        w1_rom[2630] = 2'b00;
        w1_rom[2631] = 2'b00;
        w1_rom[2632] = 2'b00;
        w1_rom[2633] = 2'b11;
        w1_rom[2634] = 2'b11;
        w1_rom[2635] = 2'b11;
        w1_rom[2636] = 2'b11;
        w1_rom[2637] = 2'b11;
        w1_rom[2638] = 2'b01;
        w1_rom[2639] = 2'b01;
        // Weights 2640-2655
        w1_rom[2640] = 2'b00;
        w1_rom[2641] = 2'b00;
        w1_rom[2642] = 2'b01;
        w1_rom[2643] = 2'b00;
        w1_rom[2644] = 2'b00;
        w1_rom[2645] = 2'b00;
        w1_rom[2646] = 2'b00;
        w1_rom[2647] = 2'b01;
        w1_rom[2648] = 2'b01;
        w1_rom[2649] = 2'b01;
        w1_rom[2650] = 2'b01;
        w1_rom[2651] = 2'b01;
        w1_rom[2652] = 2'b01;
        w1_rom[2653] = 2'b11;
        w1_rom[2654] = 2'b11;
        w1_rom[2655] = 2'b01;
        // Weights 2656-2671
        w1_rom[2656] = 2'b00;
        w1_rom[2657] = 2'b11;
        w1_rom[2658] = 2'b11;
        w1_rom[2659] = 2'b11;
        w1_rom[2660] = 2'b00;
        w1_rom[2661] = 2'b00;
        w1_rom[2662] = 2'b01;
        w1_rom[2663] = 2'b00;
        w1_rom[2664] = 2'b11;
        w1_rom[2665] = 2'b00;
        w1_rom[2666] = 2'b11;
        w1_rom[2667] = 2'b00;
        w1_rom[2668] = 2'b00;
        w1_rom[2669] = 2'b11;
        w1_rom[2670] = 2'b00;
        w1_rom[2671] = 2'b11;
        // Weights 2672-2687
        w1_rom[2672] = 2'b00;
        w1_rom[2673] = 2'b00;
        w1_rom[2674] = 2'b01;
        w1_rom[2675] = 2'b00;
        w1_rom[2676] = 2'b00;
        w1_rom[2677] = 2'b11;
        w1_rom[2678] = 2'b00;
        w1_rom[2679] = 2'b00;
        w1_rom[2680] = 2'b00;
        w1_rom[2681] = 2'b01;
        w1_rom[2682] = 2'b00;
        w1_rom[2683] = 2'b00;
        w1_rom[2684] = 2'b00;
        w1_rom[2685] = 2'b00;
        w1_rom[2686] = 2'b11;
        w1_rom[2687] = 2'b00;
        // Weights 2688-2703
        w1_rom[2688] = 2'b01;
        w1_rom[2689] = 2'b00;
        w1_rom[2690] = 2'b00;
        w1_rom[2691] = 2'b01;
        w1_rom[2692] = 2'b01;
        w1_rom[2693] = 2'b01;
        w1_rom[2694] = 2'b01;
        w1_rom[2695] = 2'b00;
        w1_rom[2696] = 2'b00;
        w1_rom[2697] = 2'b01;
        w1_rom[2698] = 2'b11;
        w1_rom[2699] = 2'b11;
        w1_rom[2700] = 2'b11;
        w1_rom[2701] = 2'b11;
        w1_rom[2702] = 2'b11;
        w1_rom[2703] = 2'b11;
        // Weights 2704-2719
        w1_rom[2704] = 2'b01;
        w1_rom[2705] = 2'b01;
        w1_rom[2706] = 2'b11;
        w1_rom[2707] = 2'b11;
        w1_rom[2708] = 2'b01;
        w1_rom[2709] = 2'b00;
        w1_rom[2710] = 2'b11;
        w1_rom[2711] = 2'b11;
        w1_rom[2712] = 2'b01;
        w1_rom[2713] = 2'b01;
        w1_rom[2714] = 2'b01;
        w1_rom[2715] = 2'b11;
        w1_rom[2716] = 2'b11;
        w1_rom[2717] = 2'b01;
        w1_rom[2718] = 2'b01;
        w1_rom[2719] = 2'b11;
        // Weights 2720-2735
        w1_rom[2720] = 2'b00;
        w1_rom[2721] = 2'b01;
        w1_rom[2722] = 2'b01;
        w1_rom[2723] = 2'b11;
        w1_rom[2724] = 2'b11;
        w1_rom[2725] = 2'b01;
        w1_rom[2726] = 2'b01;
        w1_rom[2727] = 2'b01;
        w1_rom[2728] = 2'b11;
        w1_rom[2729] = 2'b11;
        w1_rom[2730] = 2'b11;
        w1_rom[2731] = 2'b01;
        w1_rom[2732] = 2'b01;
        w1_rom[2733] = 2'b11;
        w1_rom[2734] = 2'b11;
        w1_rom[2735] = 2'b01;
        // Weights 2736-2751
        w1_rom[2736] = 2'b00;
        w1_rom[2737] = 2'b11;
        w1_rom[2738] = 2'b11;
        w1_rom[2739] = 2'b11;
        w1_rom[2740] = 2'b11;
        w1_rom[2741] = 2'b11;
        w1_rom[2742] = 2'b11;
        w1_rom[2743] = 2'b00;
        w1_rom[2744] = 2'b11;
        w1_rom[2745] = 2'b00;
        w1_rom[2746] = 2'b00;
        w1_rom[2747] = 2'b11;
        w1_rom[2748] = 2'b11;
        w1_rom[2749] = 2'b11;
        w1_rom[2750] = 2'b00;
        w1_rom[2751] = 2'b00;
        // Weights 2752-2767
        w1_rom[2752] = 2'b00;
        w1_rom[2753] = 2'b01;
        w1_rom[2754] = 2'b01;
        w1_rom[2755] = 2'b01;
        w1_rom[2756] = 2'b01;
        w1_rom[2757] = 2'b01;
        w1_rom[2758] = 2'b01;
        w1_rom[2759] = 2'b00;
        w1_rom[2760] = 2'b00;
        w1_rom[2761] = 2'b01;
        w1_rom[2762] = 2'b01;
        w1_rom[2763] = 2'b01;
        w1_rom[2764] = 2'b01;
        w1_rom[2765] = 2'b00;
        w1_rom[2766] = 2'b11;
        w1_rom[2767] = 2'b00;
        // Weights 2768-2783
        w1_rom[2768] = 2'b00;
        w1_rom[2769] = 2'b01;
        w1_rom[2770] = 2'b01;
        w1_rom[2771] = 2'b11;
        w1_rom[2772] = 2'b11;
        w1_rom[2773] = 2'b11;
        w1_rom[2774] = 2'b11;
        w1_rom[2775] = 2'b11;
        w1_rom[2776] = 2'b00;
        w1_rom[2777] = 2'b11;
        w1_rom[2778] = 2'b11;
        w1_rom[2779] = 2'b11;
        w1_rom[2780] = 2'b01;
        w1_rom[2781] = 2'b11;
        w1_rom[2782] = 2'b11;
        w1_rom[2783] = 2'b00;
        // Weights 2784-2799
        w1_rom[2784] = 2'b00;
        w1_rom[2785] = 2'b11;
        w1_rom[2786] = 2'b11;
        w1_rom[2787] = 2'b00;
        w1_rom[2788] = 2'b01;
        w1_rom[2789] = 2'b00;
        w1_rom[2790] = 2'b01;
        w1_rom[2791] = 2'b01;
        w1_rom[2792] = 2'b00;
        w1_rom[2793] = 2'b01;
        w1_rom[2794] = 2'b11;
        w1_rom[2795] = 2'b01;
        w1_rom[2796] = 2'b01;
        w1_rom[2797] = 2'b01;
        w1_rom[2798] = 2'b01;
        w1_rom[2799] = 2'b01;
        // Weights 2800-2815
        w1_rom[2800] = 2'b00;
        w1_rom[2801] = 2'b01;
        w1_rom[2802] = 2'b00;
        w1_rom[2803] = 2'b11;
        w1_rom[2804] = 2'b00;
        w1_rom[2805] = 2'b00;
        w1_rom[2806] = 2'b11;
        w1_rom[2807] = 2'b00;
        w1_rom[2808] = 2'b00;
        w1_rom[2809] = 2'b00;
        w1_rom[2810] = 2'b00;
        w1_rom[2811] = 2'b11;
        w1_rom[2812] = 2'b11;
        w1_rom[2813] = 2'b11;
        w1_rom[2814] = 2'b11;
        w1_rom[2815] = 2'b00;

        // Weights 2816-2831
        w1_rom[2816] = 2'b00;
        w1_rom[2817] = 2'b01;
        w1_rom[2818] = 2'b00;
        w1_rom[2819] = 2'b00;
        w1_rom[2820] = 2'b01;
        w1_rom[2821] = 2'b01;
        w1_rom[2822] = 2'b00;
        w1_rom[2823] = 2'b00;
        w1_rom[2824] = 2'b01;
        w1_rom[2825] = 2'b11;
        w1_rom[2826] = 2'b11;
        w1_rom[2827] = 2'b11;
        w1_rom[2828] = 2'b11;
        w1_rom[2829] = 2'b01;
        w1_rom[2830] = 2'b01;
        w1_rom[2831] = 2'b01;
        // Weights 2832-2847
        w1_rom[2832] = 2'b00;
        w1_rom[2833] = 2'b11;
        w1_rom[2834] = 2'b11;
        w1_rom[2835] = 2'b01;
        w1_rom[2836] = 2'b01;
        w1_rom[2837] = 2'b11;
        w1_rom[2838] = 2'b00;
        w1_rom[2839] = 2'b01;
        w1_rom[2840] = 2'b00;
        w1_rom[2841] = 2'b01;
        w1_rom[2842] = 2'b01;
        w1_rom[2843] = 2'b01;
        w1_rom[2844] = 2'b11;
        w1_rom[2845] = 2'b11;
        w1_rom[2846] = 2'b01;
        w1_rom[2847] = 2'b01;
        // Weights 2848-2863
        w1_rom[2848] = 2'b00;
        w1_rom[2849] = 2'b01;
        w1_rom[2850] = 2'b01;
        w1_rom[2851] = 2'b11;
        w1_rom[2852] = 2'b11;
        w1_rom[2853] = 2'b11;
        w1_rom[2854] = 2'b01;
        w1_rom[2855] = 2'b00;
        w1_rom[2856] = 2'b00;
        w1_rom[2857] = 2'b11;
        w1_rom[2858] = 2'b00;
        w1_rom[2859] = 2'b00;
        w1_rom[2860] = 2'b11;
        w1_rom[2861] = 2'b11;
        w1_rom[2862] = 2'b11;
        w1_rom[2863] = 2'b11;
        // Weights 2864-2879
        w1_rom[2864] = 2'b00;
        w1_rom[2865] = 2'b11;
        w1_rom[2866] = 2'b11;
        w1_rom[2867] = 2'b01;
        w1_rom[2868] = 2'b00;
        w1_rom[2869] = 2'b11;
        w1_rom[2870] = 2'b11;
        w1_rom[2871] = 2'b01;
        w1_rom[2872] = 2'b00;
        w1_rom[2873] = 2'b00;
        w1_rom[2874] = 2'b00;
        w1_rom[2875] = 2'b11;
        w1_rom[2876] = 2'b00;
        w1_rom[2877] = 2'b01;
        w1_rom[2878] = 2'b00;
        w1_rom[2879] = 2'b00;
        // Weights 2880-2895
        w1_rom[2880] = 2'b00;
        w1_rom[2881] = 2'b11;
        w1_rom[2882] = 2'b00;
        w1_rom[2883] = 2'b00;
        w1_rom[2884] = 2'b01;
        w1_rom[2885] = 2'b00;
        w1_rom[2886] = 2'b01;
        w1_rom[2887] = 2'b11;
        w1_rom[2888] = 2'b01;
        w1_rom[2889] = 2'b01;
        w1_rom[2890] = 2'b01;
        w1_rom[2891] = 2'b01;
        w1_rom[2892] = 2'b00;
        w1_rom[2893] = 2'b11;
        w1_rom[2894] = 2'b11;
        w1_rom[2895] = 2'b11;
        // Weights 2896-2911
        w1_rom[2896] = 2'b00;
        w1_rom[2897] = 2'b01;
        w1_rom[2898] = 2'b01;
        w1_rom[2899] = 2'b11;
        w1_rom[2900] = 2'b01;
        w1_rom[2901] = 2'b01;
        w1_rom[2902] = 2'b11;
        w1_rom[2903] = 2'b11;
        w1_rom[2904] = 2'b01;
        w1_rom[2905] = 2'b00;
        w1_rom[2906] = 2'b11;
        w1_rom[2907] = 2'b11;
        w1_rom[2908] = 2'b01;
        w1_rom[2909] = 2'b01;
        w1_rom[2910] = 2'b11;
        w1_rom[2911] = 2'b00;
        // Weights 2912-2927
        w1_rom[2912] = 2'b00;
        w1_rom[2913] = 2'b11;
        w1_rom[2914] = 2'b11;
        w1_rom[2915] = 2'b11;
        w1_rom[2916] = 2'b00;
        w1_rom[2917] = 2'b01;
        w1_rom[2918] = 2'b01;
        w1_rom[2919] = 2'b00;
        w1_rom[2920] = 2'b00;
        w1_rom[2921] = 2'b01;
        w1_rom[2922] = 2'b11;
        w1_rom[2923] = 2'b11;
        w1_rom[2924] = 2'b11;
        w1_rom[2925] = 2'b01;
        w1_rom[2926] = 2'b11;
        w1_rom[2927] = 2'b11;
        // Weights 2928-2943
        w1_rom[2928] = 2'b00;
        w1_rom[2929] = 2'b01;
        w1_rom[2930] = 2'b00;
        w1_rom[2931] = 2'b11;
        w1_rom[2932] = 2'b00;
        w1_rom[2933] = 2'b11;
        w1_rom[2934] = 2'b11;
        w1_rom[2935] = 2'b11;
        w1_rom[2936] = 2'b11;
        w1_rom[2937] = 2'b01;
        w1_rom[2938] = 2'b01;
        w1_rom[2939] = 2'b01;
        w1_rom[2940] = 2'b01;
        w1_rom[2941] = 2'b01;
        w1_rom[2942] = 2'b00;
        w1_rom[2943] = 2'b00;
        // Weights 2944-2959
        w1_rom[2944] = 2'b00;
        w1_rom[2945] = 2'b00;
        w1_rom[2946] = 2'b00;
        w1_rom[2947] = 2'b00;
        w1_rom[2948] = 2'b00;
        w1_rom[2949] = 2'b00;
        w1_rom[2950] = 2'b00;
        w1_rom[2951] = 2'b00;
        w1_rom[2952] = 2'b01;
        w1_rom[2953] = 2'b11;
        w1_rom[2954] = 2'b11;
        w1_rom[2955] = 2'b00;
        w1_rom[2956] = 2'b00;
        w1_rom[2957] = 2'b00;
        w1_rom[2958] = 2'b00;
        w1_rom[2959] = 2'b01;
        // Weights 2960-2975
        w1_rom[2960] = 2'b01;
        w1_rom[2961] = 2'b11;
        w1_rom[2962] = 2'b11;
        w1_rom[2963] = 2'b00;
        w1_rom[2964] = 2'b01;
        w1_rom[2965] = 2'b00;
        w1_rom[2966] = 2'b11;
        w1_rom[2967] = 2'b01;
        w1_rom[2968] = 2'b11;
        w1_rom[2969] = 2'b01;
        w1_rom[2970] = 2'b01;
        w1_rom[2971] = 2'b01;
        w1_rom[2972] = 2'b11;
        w1_rom[2973] = 2'b11;
        w1_rom[2974] = 2'b11;
        w1_rom[2975] = 2'b00;
        // Weights 2976-2991
        w1_rom[2976] = 2'b00;
        w1_rom[2977] = 2'b11;
        w1_rom[2978] = 2'b00;
        w1_rom[2979] = 2'b00;
        w1_rom[2980] = 2'b00;
        w1_rom[2981] = 2'b11;
        w1_rom[2982] = 2'b11;
        w1_rom[2983] = 2'b00;
        w1_rom[2984] = 2'b00;
        w1_rom[2985] = 2'b01;
        w1_rom[2986] = 2'b00;
        w1_rom[2987] = 2'b11;
        w1_rom[2988] = 2'b00;
        w1_rom[2989] = 2'b00;
        w1_rom[2990] = 2'b00;
        w1_rom[2991] = 2'b11;
        // Weights 2992-3007
        w1_rom[2992] = 2'b00;
        w1_rom[2993] = 2'b00;
        w1_rom[2994] = 2'b00;
        w1_rom[2995] = 2'b11;
        w1_rom[2996] = 2'b11;
        w1_rom[2997] = 2'b11;
        w1_rom[2998] = 2'b01;
        w1_rom[2999] = 2'b00;
        w1_rom[3000] = 2'b00;
        w1_rom[3001] = 2'b00;
        w1_rom[3002] = 2'b00;
        w1_rom[3003] = 2'b00;
        w1_rom[3004] = 2'b11;
        w1_rom[3005] = 2'b01;
        w1_rom[3006] = 2'b01;
        w1_rom[3007] = 2'b00;
        // Weights 3008-3023
        w1_rom[3008] = 2'b01;
        w1_rom[3009] = 2'b00;
        w1_rom[3010] = 2'b01;
        w1_rom[3011] = 2'b01;
        w1_rom[3012] = 2'b01;
        w1_rom[3013] = 2'b01;
        w1_rom[3014] = 2'b00;
        w1_rom[3015] = 2'b00;
        w1_rom[3016] = 2'b00;
        w1_rom[3017] = 2'b11;
        w1_rom[3018] = 2'b00;
        w1_rom[3019] = 2'b00;
        w1_rom[3020] = 2'b01;
        w1_rom[3021] = 2'b01;
        w1_rom[3022] = 2'b00;
        w1_rom[3023] = 2'b00;
        // Weights 3024-3039
        w1_rom[3024] = 2'b00;
        w1_rom[3025] = 2'b11;
        w1_rom[3026] = 2'b11;
        w1_rom[3027] = 2'b11;
        w1_rom[3028] = 2'b11;
        w1_rom[3029] = 2'b11;
        w1_rom[3030] = 2'b11;
        w1_rom[3031] = 2'b11;
        w1_rom[3032] = 2'b11;
        w1_rom[3033] = 2'b11;
        w1_rom[3034] = 2'b11;
        w1_rom[3035] = 2'b11;
        w1_rom[3036] = 2'b11;
        w1_rom[3037] = 2'b11;
        w1_rom[3038] = 2'b01;
        w1_rom[3039] = 2'b01;
        // Weights 3040-3055
        w1_rom[3040] = 2'b00;
        w1_rom[3041] = 2'b01;
        w1_rom[3042] = 2'b01;
        w1_rom[3043] = 2'b01;
        w1_rom[3044] = 2'b11;
        w1_rom[3045] = 2'b11;
        w1_rom[3046] = 2'b01;
        w1_rom[3047] = 2'b01;
        w1_rom[3048] = 2'b11;
        w1_rom[3049] = 2'b01;
        w1_rom[3050] = 2'b01;
        w1_rom[3051] = 2'b01;
        w1_rom[3052] = 2'b01;
        w1_rom[3053] = 2'b01;
        w1_rom[3054] = 2'b01;
        w1_rom[3055] = 2'b01;
        // Weights 3056-3071
        w1_rom[3056] = 2'b00;
        w1_rom[3057] = 2'b00;
        w1_rom[3058] = 2'b00;
        w1_rom[3059] = 2'b01;
        w1_rom[3060] = 2'b01;
        w1_rom[3061] = 2'b01;
        w1_rom[3062] = 2'b00;
        w1_rom[3063] = 2'b00;
        w1_rom[3064] = 2'b00;
        w1_rom[3065] = 2'b11;
        w1_rom[3066] = 2'b11;
        w1_rom[3067] = 2'b11;
        w1_rom[3068] = 2'b11;
        w1_rom[3069] = 2'b11;
        w1_rom[3070] = 2'b11;
        w1_rom[3071] = 2'b00;


        // Biases (48 entries)
        b1_rom[ 0] = 4'h2;
        b1_rom[ 1] = 4'h0;
        b1_rom[ 2] = 4'hF;
        b1_rom[ 3] = 4'h3;
        b1_rom[ 4] = 4'h4;
        b1_rom[ 5] = 4'h3;
        b1_rom[ 6] = 4'h1;
        b1_rom[ 7] = 4'h0;
        b1_rom[ 8] = 4'hC;
        b1_rom[ 9] = 4'hF;
        b1_rom[10] = 4'h0;
        b1_rom[11] = 4'h3;
        b1_rom[12] = 4'h3;
        b1_rom[13] = 4'h0;
        b1_rom[14] = 4'h0;
        b1_rom[15] = 4'h2;
        b1_rom[16] = 4'h1;
        b1_rom[17] = 4'h4;
        b1_rom[18] = 4'hB;
        b1_rom[19] = 4'h5;
        b1_rom[20] = 4'h2;
        b1_rom[21] = 4'h4;
        b1_rom[22] = 4'hD;
        b1_rom[23] = 4'h0;
        b1_rom[24] = 4'hE;
        b1_rom[25] = 4'hF;
        b1_rom[26] = 4'hF;
        b1_rom[27] = 4'h0;
        b1_rom[28] = 4'h2;
        b1_rom[29] = 4'h0;
        b1_rom[30] = 4'hF;
        b1_rom[31] = 4'h1;
        b1_rom[32] = 4'h0;
        b1_rom[33] = 4'hF;
        b1_rom[34] = 4'h1;
        b1_rom[35] = 4'h5;
        b1_rom[36] = 4'h3;
        b1_rom[37] = 4'h1;
        b1_rom[38] = 4'h1;
        b1_rom[39] = 4'h2;
        b1_rom[40] = 4'h1;
        b1_rom[41] = 4'h3;
        b1_rom[42] = 4'h7;
        b1_rom[43] = 4'h2;
        b1_rom[44] = 4'h3;
        b1_rom[45] = 4'h0;
        b1_rom[46] = 4'h3;
        b1_rom[47] = 4'h1;

    end
    
    // ========================================================================
    // FSM States
    // ========================================================================
    localparam IDLE    = 2'b00;
    localparam COMPUTE = 2'b01;
    localparam STORE   = 2'b10;
    localparam DONE_ST = 2'b11;

    reg [1:0] state;
    reg [5:0] neuron_idx;              // Current neuron (0-47)
    
    // ========================================================================
    // Output Storage
    // ========================================================================
    // Store 48 activated outputs: 48 × 2 bits = 96 bits
    reg signed [1:0] output_mem [0:47];
    
    // Output read interface - combinational
    assign read_data = output_mem[read_addr];
    
    // ========================================================================
    // Neuron Computation
    // ========================================================================
    reg neuron_start;
    wire neuron_done;
    wire signed [6:0] neuron_result;
    wire [5:0] neuron_mac_count;       // Which MAC the neuron is on
    
    // ROM addressing for current neuron - use neuron's counter
    wire [11:0] weight_addr = neuron_idx * 12'd64 + {6'd0, neuron_mac_count};
    wire [1:0] current_weight = w1_rom[weight_addr];
    wire signed [3:0] current_bias = $signed(b1_rom[neuron_idx]);
    
    // Read pixel directly from array using neuron's MAC count
    wire [1:0] current_pixel = pixels[neuron_mac_count];
    
    layer1_neuron neuron (
        .clk(clk),
        .rst_n(rst_n),
        .start(neuron_start),
        .input_val(current_pixel),       // Read directly from pixel array
        .weight(current_weight),
        .bias(current_bias),
        .done(neuron_done),
        .result(neuron_result),
        .mac_count_out(neuron_mac_count) // Get neuron's MAC counter
    );
    
    // ========================================================================
    // Activation
    // ========================================================================
    wire signed [1:0] activated_result;
    
    sign_activation activation (
        .in_val(neuron_result),
        .out(activated_result)
    );
    
    // ========================================================================
    // FSM and Control
    // ========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            neuron_idx <= 6'd0;
            neuron_start <= 1'b0;
            done <= 1'b0;
            busy <= 1'b0;
        end else begin
            case (state)
                IDLE: begin
                    done <= 1'b0;
                    busy <= 1'b0;
                    neuron_start <= 1'b0;
                    
                    if (start) begin
                        neuron_idx <= 6'd0;
                        state <= COMPUTE;
                        neuron_start <= 1'b1;  // Start first neuron
                        busy <= 1'b1;
                    end
                end
                
                COMPUTE: begin
                    neuron_start <= 1'b0;  // Clear start after one cycle
                    
                    // No counter management needed - neuron tracks its own MAC count!
                    
                    if (neuron_done) begin
                        // Store activated result
                        output_mem[neuron_idx] <= activated_result;
                        state <= STORE;
                    end
                end
                
                STORE: begin
                    // Check if more neurons to process
                    if (neuron_idx < 6'd47) begin
                        neuron_idx <= neuron_idx + 1'b1;
                        state <= COMPUTE;
                        neuron_start <= 1'b1;  // Start next neuron
                    end else begin
                        // All neurons done
                        state <= DONE_ST;
                        done <= 1'b1;
                        busy <= 1'b0;
                    end
                end
                
                DONE_ST: begin
                    // Stay in DONE until start goes low
                    if (!start) begin
                        state <= IDLE;
                    end
                end
                
                default: state <= IDLE;
            endcase
        end
    end

endmodule
