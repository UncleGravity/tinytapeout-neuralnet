/*
 * Layer 2 Full - Complete second layer with integrated ROM
 * 
 * Self-contained module that processes all 10 output neurons sequentially.
 * Weights and biases are stored in internal ROM (loaded from hex files).
 * 
 * Input: 48 signed activations from Layer 1 (streamed cyclically by parent)
 * Output: 10 signed 6-bit logits stored internally, readable after done
 * 
 * Architecture:
 *   - Internal ROM: W2 weights (480 entries) + b2 biases (10 entries)
 *   - Reuses 1 layer2_neuron for all 10 outputs
 *   - FSM manages sequential processing and ROM addressing
 * 
 * Memory:
 *   - W2: 480 weights × 2 bits = 960 bits
 *   - b2: 10 biases × 4 bits = 40 bits
 *   - Output buffer: 10 × 6 bits = 60 bits
 *   - Total: 1,060 bits (133 bytes)
 * 
 * Timing:
 *   - Each neuron: ~52 cycles (48 MACs + bias + overhead)
 *   - Total: ~520 cycles for all 10 neurons
 */

module layer2_full (
    input  wire        clk,
    input  wire        rst_n,
    input  wire        start,              // Start Layer 2 computation
    input  wire [95:0] layer1_activations_flat, // All 48 Layer 1 outputs as flat vector (48 × 2-bit = 96 bits)
    output reg         done,               // Computation complete
    output reg         busy,               // Currently computing
    // Read interface for outputs (after done=1)
    input  wire [3:0]  read_addr,          // Which output to read (0-9)
    output wire signed [5:0] read_data     // Logit value at read_addr
);

    // ========================================================================
    // Unpack flat activation vector into array
    // ========================================================================
    reg signed [1:0] layer1_activations [0:47];
    integer k;
    always @(*) begin
        for (k = 0; k < 48; k = k + 1) begin
            layer1_activations[k] = layer1_activations_flat[k*2 +: 2];
        end
    end

    // ========================================================================
    // Weight and Bias ROM
    // ========================================================================
    
    // Layer 2 Weight ROM: 480 weights (10 neurons × 48 inputs)
    // Column-major: neuron N weights at addresses [N*48, N*48+47]
    reg [1:0] w2_rom [0:479];
    
    // Layer 2 Bias ROM: 10 biases
    reg [3:0] b2_rom [0:9];
    
    // Inline initialization - generated from weights.npz
    // This works for both RTL and gate-level simulation
    initial begin
        // Weights (480 entries: 10 neurons × 48 inputs)
        // Weights   0- 15
        w2_rom[  0] = 2'b00;
        w2_rom[  1] = 2'b11;
        w2_rom[  2] = 2'b00;
        w2_rom[  3] = 2'b11;
        w2_rom[  4] = 2'b00;
        w2_rom[  5] = 2'b11;
        w2_rom[  6] = 2'b00;
        w2_rom[  7] = 2'b00;
        w2_rom[  8] = 2'b11;
        w2_rom[  9] = 2'b00;
        w2_rom[ 10] = 2'b00;
        w2_rom[ 11] = 2'b00;
        w2_rom[ 12] = 2'b11;
        w2_rom[ 13] = 2'b00;
        w2_rom[ 14] = 2'b11;
        w2_rom[ 15] = 2'b11;
        // Weights  16- 31
        w2_rom[ 16] = 2'b01;
        w2_rom[ 17] = 2'b00;
        w2_rom[ 18] = 2'b11;
        w2_rom[ 19] = 2'b00;
        w2_rom[ 20] = 2'b00;
        w2_rom[ 21] = 2'b00;
        w2_rom[ 22] = 2'b00;
        w2_rom[ 23] = 2'b00;
        w2_rom[ 24] = 2'b01;
        w2_rom[ 25] = 2'b00;
        w2_rom[ 26] = 2'b11;
        w2_rom[ 27] = 2'b11;
        w2_rom[ 28] = 2'b00;
        w2_rom[ 29] = 2'b00;
        w2_rom[ 30] = 2'b00;
        w2_rom[ 31] = 2'b00;
        // Weights  32- 47
        w2_rom[ 32] = 2'b00;
        w2_rom[ 33] = 2'b00;
        w2_rom[ 34] = 2'b01;
        w2_rom[ 35] = 2'b00;
        w2_rom[ 36] = 2'b00;
        w2_rom[ 37] = 2'b00;
        w2_rom[ 38] = 2'b00;
        w2_rom[ 39] = 2'b00;
        w2_rom[ 40] = 2'b00;
        w2_rom[ 41] = 2'b00;
        w2_rom[ 42] = 2'b00;
        w2_rom[ 43] = 2'b11;
        w2_rom[ 44] = 2'b01;
        w2_rom[ 45] = 2'b00;
        w2_rom[ 46] = 2'b00;
        w2_rom[ 47] = 2'b01;
        // Weights  48- 63
        w2_rom[ 48] = 2'b00;
        w2_rom[ 49] = 2'b01;
        w2_rom[ 50] = 2'b00;
        w2_rom[ 51] = 2'b11;
        w2_rom[ 52] = 2'b01;
        w2_rom[ 53] = 2'b00;
        w2_rom[ 54] = 2'b00;
        w2_rom[ 55] = 2'b11;
        w2_rom[ 56] = 2'b00;
        w2_rom[ 57] = 2'b00;
        w2_rom[ 58] = 2'b00;
        w2_rom[ 59] = 2'b00;
        w2_rom[ 60] = 2'b01;
        w2_rom[ 61] = 2'b00;
        w2_rom[ 62] = 2'b00;
        w2_rom[ 63] = 2'b11;
        // Weights  64- 79
        w2_rom[ 64] = 2'b00;
        w2_rom[ 65] = 2'b00;
        w2_rom[ 66] = 2'b00;
        w2_rom[ 67] = 2'b00;
        w2_rom[ 68] = 2'b01;
        w2_rom[ 69] = 2'b01;
        w2_rom[ 70] = 2'b11;
        w2_rom[ 71] = 2'b11;
        w2_rom[ 72] = 2'b11;
        w2_rom[ 73] = 2'b00;
        w2_rom[ 74] = 2'b01;
        w2_rom[ 75] = 2'b01;
        w2_rom[ 76] = 2'b00;
        w2_rom[ 77] = 2'b00;
        w2_rom[ 78] = 2'b00;
        w2_rom[ 79] = 2'b00;
        // Weights  80- 95
        w2_rom[ 80] = 2'b00;
        w2_rom[ 81] = 2'b00;
        w2_rom[ 82] = 2'b11;
        w2_rom[ 83] = 2'b00;
        w2_rom[ 84] = 2'b00;
        w2_rom[ 85] = 2'b00;
        w2_rom[ 86] = 2'b00;
        w2_rom[ 87] = 2'b00;
        w2_rom[ 88] = 2'b00;
        w2_rom[ 89] = 2'b01;
        w2_rom[ 90] = 2'b00;
        w2_rom[ 91] = 2'b01;
        w2_rom[ 92] = 2'b00;
        w2_rom[ 93] = 2'b00;
        w2_rom[ 94] = 2'b00;
        w2_rom[ 95] = 2'b00;
        // Weights  96-111
        w2_rom[ 96] = 2'b01;
        w2_rom[ 97] = 2'b00;
        w2_rom[ 98] = 2'b00;
        w2_rom[ 99] = 2'b00;
        w2_rom[100] = 2'b00;
        w2_rom[101] = 2'b01;
        w2_rom[102] = 2'b00;
        w2_rom[103] = 2'b11;
        w2_rom[104] = 2'b00;
        w2_rom[105] = 2'b11;
        w2_rom[106] = 2'b00;
        w2_rom[107] = 2'b00;
        w2_rom[108] = 2'b01;
        w2_rom[109] = 2'b00;
        w2_rom[110] = 2'b11;
        w2_rom[111] = 2'b00;
        // Weights 112-127
        w2_rom[112] = 2'b00;
        w2_rom[113] = 2'b00;
        w2_rom[114] = 2'b01;
        w2_rom[115] = 2'b00;
        w2_rom[116] = 2'b01;
        w2_rom[117] = 2'b01;
        w2_rom[118] = 2'b00;
        w2_rom[119] = 2'b00;
        w2_rom[120] = 2'b01;
        w2_rom[121] = 2'b00;
        w2_rom[122] = 2'b00;
        w2_rom[123] = 2'b11;
        w2_rom[124] = 2'b00;
        w2_rom[125] = 2'b01;
        w2_rom[126] = 2'b00;
        w2_rom[127] = 2'b00;

        // Weights 128-143
        w2_rom[128] = 2'b00;
        w2_rom[129] = 2'b00;
        w2_rom[130] = 2'b00;
        w2_rom[131] = 2'b11;
        w2_rom[132] = 2'b00;
        w2_rom[133] = 2'b00;
        w2_rom[134] = 2'b00;
        w2_rom[135] = 2'b00;
        w2_rom[136] = 2'b00;
        w2_rom[137] = 2'b00;
        w2_rom[138] = 2'b00;
        w2_rom[139] = 2'b01;
        w2_rom[140] = 2'b11;
        w2_rom[141] = 2'b01;
        w2_rom[142] = 2'b00;
        w2_rom[143] = 2'b00;
        // Weights 144-159
        w2_rom[144] = 2'b01;
        w2_rom[145] = 2'b00;
        w2_rom[146] = 2'b00;
        w2_rom[147] = 2'b11;
        w2_rom[148] = 2'b00;
        w2_rom[149] = 2'b00;
        w2_rom[150] = 2'b00;
        w2_rom[151] = 2'b00;
        w2_rom[152] = 2'b00;
        w2_rom[153] = 2'b00;
        w2_rom[154] = 2'b01;
        w2_rom[155] = 2'b00;
        w2_rom[156] = 2'b01;
        w2_rom[157] = 2'b00;
        w2_rom[158] = 2'b00;
        w2_rom[159] = 2'b11;
        // Weights 160-175
        w2_rom[160] = 2'b00;
        w2_rom[161] = 2'b01;
        w2_rom[162] = 2'b00;
        w2_rom[163] = 2'b00;
        w2_rom[164] = 2'b00;
        w2_rom[165] = 2'b00;
        w2_rom[166] = 2'b00;
        w2_rom[167] = 2'b11;
        w2_rom[168] = 2'b01;
        w2_rom[169] = 2'b00;
        w2_rom[170] = 2'b11;
        w2_rom[171] = 2'b00;
        w2_rom[172] = 2'b00;
        w2_rom[173] = 2'b00;
        w2_rom[174] = 2'b00;
        w2_rom[175] = 2'b00;
        // Weights 176-191
        w2_rom[176] = 2'b00;
        w2_rom[177] = 2'b00;
        w2_rom[178] = 2'b00;
        w2_rom[179] = 2'b11;
        w2_rom[180] = 2'b00;
        w2_rom[181] = 2'b01;
        w2_rom[182] = 2'b00;
        w2_rom[183] = 2'b00;
        w2_rom[184] = 2'b00;
        w2_rom[185] = 2'b00;
        w2_rom[186] = 2'b11;
        w2_rom[187] = 2'b01;
        w2_rom[188] = 2'b11;
        w2_rom[189] = 2'b01;
        w2_rom[190] = 2'b00;
        w2_rom[191] = 2'b11;
        // Weights 192-207
        w2_rom[192] = 2'b00;
        w2_rom[193] = 2'b00;
        w2_rom[194] = 2'b00;
        w2_rom[195] = 2'b01;
        w2_rom[196] = 2'b00;
        w2_rom[197] = 2'b01;
        w2_rom[198] = 2'b00;
        w2_rom[199] = 2'b00;
        w2_rom[200] = 2'b01;
        w2_rom[201] = 2'b00;
        w2_rom[202] = 2'b00;
        w2_rom[203] = 2'b01;
        w2_rom[204] = 2'b00;
        w2_rom[205] = 2'b00;
        w2_rom[206] = 2'b00;
        w2_rom[207] = 2'b01;
        // Weights 208-223
        w2_rom[208] = 2'b01;
        w2_rom[209] = 2'b11;
        w2_rom[210] = 2'b11;
        w2_rom[211] = 2'b00;
        w2_rom[212] = 2'b01;
        w2_rom[213] = 2'b11;
        w2_rom[214] = 2'b00;
        w2_rom[215] = 2'b11;
        w2_rom[216] = 2'b11;
        w2_rom[217] = 2'b11;
        w2_rom[218] = 2'b01;
        w2_rom[219] = 2'b00;
        w2_rom[220] = 2'b00;
        w2_rom[221] = 2'b01;
        w2_rom[222] = 2'b00;
        w2_rom[223] = 2'b01;
        // Weights 224-239
        w2_rom[224] = 2'b00;
        w2_rom[225] = 2'b00;
        w2_rom[226] = 2'b00;
        w2_rom[227] = 2'b01;
        w2_rom[228] = 2'b11;
        w2_rom[229] = 2'b00;
        w2_rom[230] = 2'b00;
        w2_rom[231] = 2'b00;
        w2_rom[232] = 2'b00;
        w2_rom[233] = 2'b00;
        w2_rom[234] = 2'b01;
        w2_rom[235] = 2'b00;
        w2_rom[236] = 2'b00;
        w2_rom[237] = 2'b00;
        w2_rom[238] = 2'b00;
        w2_rom[239] = 2'b00;
        // Weights 240-255
        w2_rom[240] = 2'b00;
        w2_rom[241] = 2'b00;
        w2_rom[242] = 2'b00;
        w2_rom[243] = 2'b00;
        w2_rom[244] = 2'b00;
        w2_rom[245] = 2'b00;
        w2_rom[246] = 2'b00;
        w2_rom[247] = 2'b00;
        w2_rom[248] = 2'b01;
        w2_rom[249] = 2'b00;
        w2_rom[250] = 2'b01;
        w2_rom[251] = 2'b01;
        w2_rom[252] = 2'b00;
        w2_rom[253] = 2'b00;
        w2_rom[254] = 2'b11;
        w2_rom[255] = 2'b11;

        // Weights 256-271
        w2_rom[256] = 2'b01;
        w2_rom[257] = 2'b00;
        w2_rom[258] = 2'b00;
        w2_rom[259] = 2'b00;
        w2_rom[260] = 2'b00;
        w2_rom[261] = 2'b00;
        w2_rom[262] = 2'b00;
        w2_rom[263] = 2'b00;
        w2_rom[264] = 2'b01;
        w2_rom[265] = 2'b00;
        w2_rom[266] = 2'b01;
        w2_rom[267] = 2'b00;
        w2_rom[268] = 2'b00;
        w2_rom[269] = 2'b00;
        w2_rom[270] = 2'b00;
        w2_rom[271] = 2'b00;
        // Weights 272-287
        w2_rom[272] = 2'b00;
        w2_rom[273] = 2'b00;
        w2_rom[274] = 2'b01;
        w2_rom[275] = 2'b00;
        w2_rom[276] = 2'b00;
        w2_rom[277] = 2'b11;
        w2_rom[278] = 2'b01;
        w2_rom[279] = 2'b00;
        w2_rom[280] = 2'b00;
        w2_rom[281] = 2'b01;
        w2_rom[282] = 2'b00;
        w2_rom[283] = 2'b00;
        w2_rom[284] = 2'b00;
        w2_rom[285] = 2'b00;
        w2_rom[286] = 2'b00;
        w2_rom[287] = 2'b11;
        // Weights 288-303
        w2_rom[288] = 2'b00;
        w2_rom[289] = 2'b00;
        w2_rom[290] = 2'b00;
        w2_rom[291] = 2'b01;
        w2_rom[292] = 2'b11;
        w2_rom[293] = 2'b00;
        w2_rom[294] = 2'b00;
        w2_rom[295] = 2'b11;
        w2_rom[296] = 2'b11;
        w2_rom[297] = 2'b00;
        w2_rom[298] = 2'b11;
        w2_rom[299] = 2'b00;
        w2_rom[300] = 2'b00;
        w2_rom[301] = 2'b00;
        w2_rom[302] = 2'b00;
        w2_rom[303] = 2'b00;
        // Weights 304-319
        w2_rom[304] = 2'b00;
        w2_rom[305] = 2'b11;
        w2_rom[306] = 2'b00;
        w2_rom[307] = 2'b11;
        w2_rom[308] = 2'b01;
        w2_rom[309] = 2'b11;
        w2_rom[310] = 2'b00;
        w2_rom[311] = 2'b00;
        w2_rom[312] = 2'b11;
        w2_rom[313] = 2'b01;
        w2_rom[314] = 2'b01;
        w2_rom[315] = 2'b00;
        w2_rom[316] = 2'b00;
        w2_rom[317] = 2'b01;
        w2_rom[318] = 2'b00;
        w2_rom[319] = 2'b00;
        // Weights 320-335
        w2_rom[320] = 2'b00;
        w2_rom[321] = 2'b00;
        w2_rom[322] = 2'b01;
        w2_rom[323] = 2'b11;
        w2_rom[324] = 2'b00;
        w2_rom[325] = 2'b11;
        w2_rom[326] = 2'b01;
        w2_rom[327] = 2'b11;
        w2_rom[328] = 2'b00;
        w2_rom[329] = 2'b00;
        w2_rom[330] = 2'b01;
        w2_rom[331] = 2'b01;
        w2_rom[332] = 2'b00;
        w2_rom[333] = 2'b11;
        w2_rom[334] = 2'b00;
        w2_rom[335] = 2'b01;
        // Weights 336-351
        w2_rom[336] = 2'b00;
        w2_rom[337] = 2'b00;
        w2_rom[338] = 2'b00;
        w2_rom[339] = 2'b00;
        w2_rom[340] = 2'b01;
        w2_rom[341] = 2'b00;
        w2_rom[342] = 2'b00;
        w2_rom[343] = 2'b00;
        w2_rom[344] = 2'b00;
        w2_rom[345] = 2'b01;
        w2_rom[346] = 2'b00;
        w2_rom[347] = 2'b01;
        w2_rom[348] = 2'b11;
        w2_rom[349] = 2'b00;
        w2_rom[350] = 2'b00;
        w2_rom[351] = 2'b01;
        // Weights 352-367
        w2_rom[352] = 2'b11;
        w2_rom[353] = 2'b00;
        w2_rom[354] = 2'b00;
        w2_rom[355] = 2'b00;
        w2_rom[356] = 2'b11;
        w2_rom[357] = 2'b00;
        w2_rom[358] = 2'b00;
        w2_rom[359] = 2'b11;
        w2_rom[360] = 2'b00;
        w2_rom[361] = 2'b00;
        w2_rom[362] = 2'b11;
        w2_rom[363] = 2'b00;
        w2_rom[364] = 2'b00;
        w2_rom[365] = 2'b00;
        w2_rom[366] = 2'b00;
        w2_rom[367] = 2'b00;
        // Weights 368-383
        w2_rom[368] = 2'b00;
        w2_rom[369] = 2'b11;
        w2_rom[370] = 2'b00;
        w2_rom[371] = 2'b01;
        w2_rom[372] = 2'b01;
        w2_rom[373] = 2'b00;
        w2_rom[374] = 2'b00;
        w2_rom[375] = 2'b00;
        w2_rom[376] = 2'b00;
        w2_rom[377] = 2'b01;
        w2_rom[378] = 2'b01;
        w2_rom[379] = 2'b00;
        w2_rom[380] = 2'b00;
        w2_rom[381] = 2'b01;
        w2_rom[382] = 2'b00;
        w2_rom[383] = 2'b11;

        // Weights 384-399
        w2_rom[384] = 2'b01;
        w2_rom[385] = 2'b01;
        w2_rom[386] = 2'b00;
        w2_rom[387] = 2'b00;
        w2_rom[388] = 2'b00;
        w2_rom[389] = 2'b00;
        w2_rom[390] = 2'b00;
        w2_rom[391] = 2'b00;
        w2_rom[392] = 2'b01;
        w2_rom[393] = 2'b01;
        w2_rom[394] = 2'b00;
        w2_rom[395] = 2'b00;
        w2_rom[396] = 2'b11;
        w2_rom[397] = 2'b00;
        w2_rom[398] = 2'b11;
        w2_rom[399] = 2'b11;
        // Weights 400-415
        w2_rom[400] = 2'b00;
        w2_rom[401] = 2'b11;
        w2_rom[402] = 2'b01;
        w2_rom[403] = 2'b11;
        w2_rom[404] = 2'b00;
        w2_rom[405] = 2'b11;
        w2_rom[406] = 2'b00;
        w2_rom[407] = 2'b01;
        w2_rom[408] = 2'b01;
        w2_rom[409] = 2'b00;
        w2_rom[410] = 2'b01;
        w2_rom[411] = 2'b00;
        w2_rom[412] = 2'b00;
        w2_rom[413] = 2'b00;
        w2_rom[414] = 2'b00;
        w2_rom[415] = 2'b00;
        // Weights 416-431
        w2_rom[416] = 2'b01;
        w2_rom[417] = 2'b00;
        w2_rom[418] = 2'b00;
        w2_rom[419] = 2'b00;
        w2_rom[420] = 2'b01;
        w2_rom[421] = 2'b00;
        w2_rom[422] = 2'b00;
        w2_rom[423] = 2'b00;
        w2_rom[424] = 2'b00;
        w2_rom[425] = 2'b00;
        w2_rom[426] = 2'b11;
        w2_rom[427] = 2'b00;
        w2_rom[428] = 2'b11;
        w2_rom[429] = 2'b00;
        w2_rom[430] = 2'b00;
        w2_rom[431] = 2'b11;
        // Weights 432-447
        w2_rom[432] = 2'b00;
        w2_rom[433] = 2'b00;
        w2_rom[434] = 2'b00;
        w2_rom[435] = 2'b01;
        w2_rom[436] = 2'b01;
        w2_rom[437] = 2'b00;
        w2_rom[438] = 2'b11;
        w2_rom[439] = 2'b00;
        w2_rom[440] = 2'b01;
        w2_rom[441] = 2'b01;
        w2_rom[442] = 2'b00;
        w2_rom[443] = 2'b00;
        w2_rom[444] = 2'b00;
        w2_rom[445] = 2'b00;
        w2_rom[446] = 2'b00;
        w2_rom[447] = 2'b00;
        // Weights 448-463
        w2_rom[448] = 2'b00;
        w2_rom[449] = 2'b00;
        w2_rom[450] = 2'b00;
        w2_rom[451] = 2'b00;
        w2_rom[452] = 2'b11;
        w2_rom[453] = 2'b00;
        w2_rom[454] = 2'b00;
        w2_rom[455] = 2'b11;
        w2_rom[456] = 2'b11;
        w2_rom[457] = 2'b00;
        w2_rom[458] = 2'b00;
        w2_rom[459] = 2'b00;
        w2_rom[460] = 2'b00;
        w2_rom[461] = 2'b00;
        w2_rom[462] = 2'b00;
        w2_rom[463] = 2'b00;
        // Weights 464-479
        w2_rom[464] = 2'b00;
        w2_rom[465] = 2'b00;
        w2_rom[466] = 2'b11;
        w2_rom[467] = 2'b01;
        w2_rom[468] = 2'b00;
        w2_rom[469] = 2'b00;
        w2_rom[470] = 2'b00;
        w2_rom[471] = 2'b00;
        w2_rom[472] = 2'b00;
        w2_rom[473] = 2'b00;
        w2_rom[474] = 2'b01;
        w2_rom[475] = 2'b11;
        w2_rom[476] = 2'b00;
        w2_rom[477] = 2'b00;
        w2_rom[478] = 2'b00;
        w2_rom[479] = 2'b11;

        // Biases (10 entries)
        b2_rom[0] = 4'hE;
        b2_rom[1] = 4'hF;
        b2_rom[2] = 4'h0;
        b2_rom[3] = 4'h1;
        b2_rom[4] = 4'hF;
        b2_rom[5] = 4'h3;
        b2_rom[6] = 4'hE;
        b2_rom[7] = 4'hF;
        b2_rom[8] = 4'h2;
        b2_rom[9] = 4'h0;

    end
    
    // ========================================================================
    // FSM States
    // ========================================================================
    localparam IDLE    = 2'b00;
    localparam COMPUTE = 2'b01;
    localparam STORE   = 2'b10;
    localparam DONE_ST = 2'b11;

    reg [1:0] state;
    reg [3:0] neuron_idx;     // Current neuron (0-9)
    
    // ========================================================================
    // Output Storage
    // ========================================================================
    // Store 10 logits: 10 × 6 bits = 60 bits
    reg signed [5:0] output_mem [0:9];
    
    // Output read interface - combinational
    assign read_data = output_mem[read_addr];
    
    // ========================================================================
    // Neuron Computation
    // ========================================================================
    reg neuron_start;
    wire neuron_done;
    wire signed [5:0] neuron_result;
    wire [5:0] neuron_mac_count;  // From neuron module
    
    // ROM addressing for current neuron - use neuron's counter
    wire [8:0] weight_addr = neuron_idx * 9'd48 + {3'd0, neuron_mac_count};
    wire [1:0] current_weight = w2_rom[weight_addr];
    wire signed [3:0] current_bias = $signed(b2_rom[neuron_idx]);
    
    // Read layer1 activation directly from array using neuron's MAC count
    wire signed [1:0] current_activation = layer1_activations[neuron_mac_count];
    
    layer2_neuron neuron (
        .clk(clk),
        .rst_n(rst_n),
        .start(neuron_start),
        .input_val(current_activation),  // Read directly from layer1 array
        .weight(current_weight),
        .bias(current_bias),
        .done(neuron_done),
        .result(neuron_result),
        .mac_count_out(neuron_mac_count)
    );
    
    // ========================================================================
    // FSM and Control
    // ========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            neuron_idx <= 4'd0;
            neuron_start <= 1'b0;
            done <= 1'b0;
            busy <= 1'b0;
        end else begin
            case (state)
                IDLE: begin
                    done <= 1'b0;
                    busy <= 1'b0;
                    neuron_start <= 1'b0;
                    
                    if (start) begin
                        neuron_idx <= 4'd0;
                        state <= COMPUTE;
                        neuron_start <= 1'b1;  // Start first neuron
                        busy <= 1'b1;
                    end
                end
                
                COMPUTE: begin
                    neuron_start <= 1'b0;  // Clear start after one cycle
                    
                    // No counter management - neuron tracks its own MAC count!
                    
                    if (neuron_done) begin
                        // Store result
                        output_mem[neuron_idx] <= neuron_result;
                        state <= STORE;
                    end
                end
                
                STORE: begin
                    // Check if more neurons to process
                    if (neuron_idx < 4'd9) begin
                        neuron_idx <= neuron_idx + 1;
                        state <= COMPUTE;
                        neuron_start <= 1'b1;  // Start next neuron
                    end else begin
                        // All neurons done
                        state <= DONE_ST;
                        done <= 1'b1;
                        busy <= 1'b0;
                    end
                end
                
                DONE_ST: begin
                    // Stay in DONE until start goes low
                    if (!start) begin
                        state <= IDLE;
                    end
                end
                
                default: state <= IDLE;
            endcase
        end
    end

endmodule
